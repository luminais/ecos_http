# ====================================================================
#
#      aim711_wallclock_drivers.cdl
#
#      Wallclock drivers - support for DS1339 RTC on the 
#      ARM Industrial Module AIM 711
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002, 2003 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      rcassebohm
# Contributors:   rcassebohm
# Date:           2003-10-05
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVICES_WALLCLOCK_ARM_AIM711 {
    display       "ARM Industrial Module AIM 711 RTC Driver"
    description   "RTC driver for the ARM Industrial Module AIM 711."

    parent        CYGPKG_IO_WALLCLOCK
    active_if     CYGPKG_IO_WALLCLOCK
    active_if     CYGPKG_HAL_ARM_AIM711
    requires      CYGPKG_DEVICES_WALLCLOCK_DALLAS_DS1307

    include_dir   cyg/io

    define_proc {
        puts $::cdl_system_header "/***** AIM 711 RTC driver proc output start *****/"
        puts $::cdl_system_header "#define CYGDAT_DEVS_WALLCLOCK_DALLAS_1307_INL <cyg/io/devs_wallclock_arm_aim711.inl>"
        puts $::cdl_system_header "#define CYGDAT_DEVS_WALLCLOCK_ARM_AIM711_CFG <pkgconf/devices_wallclock_arm_aim711.h>"
        puts $::cdl_system_header "/***** AIM 711 RTC driver proc output end  *****/"
    }
}
