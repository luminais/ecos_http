# ====================================================================
#
#      flash_ea2468.cdl
#
#      FLASH memory - Hardware support on EA LPC2468 OEM board
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002, 2003 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Uwe Kindler 
# Contributors:
# Date:           2008-07-07
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_FLASH_EA2468 {
    display       "EA LPC2468 OEM board FLASH memory support"
    description   "FLASH memory device support for Embedded Artists LPC2468 OEM board"
    
    parent        CYGPKG_IO_FLASH
    active_if	  CYGPKG_IO_FLASH
    requires      CYGPKG_HAL_ARM_LPC24XX
    
    compile       -library=libextras.a flash_ea2468.c
    
    # Arguably this should do in the generic package
    # but then there is a logic loop so you can never enable it.
    cdl_interface CYGINT_DEVS_FLASH_SST_39VFXXX_REQUIRED {
        display   "Generic SST 39VFXXX driver required"
    }
    
    implements CYGINT_DEVS_FLASH_SST_39VFXXX_REQUIRED
    requires   !CYGSEM_REDBOOT_FLASH_COMBINED_FIS_AND_CONFIG
    requires   CYGNUM_REDBOOT_FLASH_CONFIG_SIZE <= 4096
    requires   {(CYGNUM_REDBOOT_FIS_DIRECTORY_ENTRY_SIZE *
                 CYGNUM_REDBOOT_FIS_DIRECTORY_ENTRY_COUNT) <= 4096}
}

# EOF flash_ea2468.cdl
