# ====================================================================
#
#      pcmcia_ipaq.cdl
#
#      PCMCIA (Compact Flash) - Hardware support on iPAQ
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      gthomas
# Original data:  gthomas
# Contributors:
#                 Richard Panton <richard.panton@3glab.com>
# Date:           2001-02-24
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_PCMCIA_IPAQ {
    display       "SA11x0/iPaq PCMCIA support"

    parent        CYGPKG_IO_PCMCIA
    active_if	  CYGPKG_IO_PCMCIA
    active_if	  CYGPKG_HAL_ARM_SA11X0_IPAQ

    implements    CYGHWR_IO_PCMCIA_DEVICE

    include_dir   .
    include_files ; # none _exported_ whatsoever
    description   "PCMCIA (Compact Flash) device support for SA11x0/iPAQ"
    compile       ipaq_pcmcia.c
}
