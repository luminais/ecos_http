# ====================================================================
#
#      ser_freescale_esci.cdl
#
#      eCos serial Freescale/esci configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002, 2006 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Ilija Koco <ilijak@siva.com.mk>
# Original data:
# Contributors:
# Date:           2006-04-20
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_IO_SERIAL_FREESCALE_ESCI {
    display       "eSCI device driver"

    parent        CYGPKG_IO_SERIAL_DEVICES
    active_if     CYGPKG_IO_SERIAL

    requires      CYGPKG_IO_SERIAL_FREESCALE_ESCI_H
    
    requires      (CYGPKG_ERROR && (CYGPKG_IO_SERIAL_FREESCALE_ESCI_A || \
                                    CYGPKG_IO_SERIAL_FREESCALE_ESCI_B || \
                                    CYGPKG_IO_SERIAL_FREESCALE_ESCI_C || \
                                    CYGPKG_IO_SERIAL_FREESCALE_ESCI_D) \
                                    )
    
    include_dir   cyg/devs

    description   "
           This option enables the serial device drivers for the
           Freescale eSCI - Enhanced Serial Communication Interface.
           eSCI is on-chip serial controller found on some freescale 
           microcontrollers such as: MAC7100 familly, etc.
           "
    compile       -library=libextras.a   ser_esci.c

    define_proc {
        puts $::cdl_system_header "/***** serial driver proc output start *****/"
        puts $::cdl_system_header "#define CYGDAT_IO_SERIAL_DEVICE_HEADER <pkgconf/io_serial_freescale_esci.h>"
        puts $::cdl_system_header "/*****  serial driver proc output end  *****/"
    }

    cdl_component CYGPKG_IO_SERIAL_FREESCALE_ESCI_A {
        display       "eSCI port A driver"
        flavor        bool
        default_value 0
        description   "
            This option includes the serial device driver for the eSCI port A."

        cdl_option CYGDAT_IO_SERIAL_FREESCALE_ESCI_A_NAME {
            display       "Device name for eSCI port A"
            flavor        data
            default_value {"\"/dev/ser0\""}
            description   "
                This option specifies the device name for the eSCI port A."
        }

        cdl_option CYGNUM_IO_SERIAL_FREESCALE_ESCI_A_BAUD {
            display       "Baud rate for the eSCI serial port A driver"
            flavor        data
            legal_values  { 300 600 1200 2400 4800 9600 14400 19200 38400 
                            57600 115200 }
            default_value 38400
            description "
                This option specifies the default baud rate (speed) for the 
                eSCI port A."
        }

        cdl_option CYGNUM_IO_SERIAL_FREESCALE_ESCI_A_BUFSIZE {
            display       "Buffer size for the sSCI port A driver"
            flavor        data
            legal_values  0 to 8192
            default_value 128
            description   "
                This option specifies the size of the internal buffers used 
                for the eSCI port A."
        }
    
        cdl_option CYGNUM_IO_SERIAL_FREESCALE_ESCI_A_INT_PRIORITY {
            display      "eSCI port A INTC priority"
            flavor       data
            legal_values 0 to 15
            default_value   7
            description "
                INTC has 16 interrupt levels: 0 (lowest) to 15 (highest).
            "
        }       
    }

    cdl_component CYGPKG_IO_SERIAL_FREESCALE_ESCI_B {
        display       "eSCI port B driver"
        flavor        bool
        default_value 0
        description   "
            This option includes the serial device driver for the eSCI port B."

        cdl_option CYGDAT_IO_SERIAL_FREESCALE_ESCI_B_NAME {
            display       "Device name for eSCI port B"
            flavor        data
            default_value {"\"/dev/ser1\""}
            description   "
                This option specifies the device name for the eSCI port B."
        }

        cdl_option CYGNUM_IO_SERIAL_FREESCALE_ESCI_B_BAUD {
            display       "Baud rate for the eSCI serial port A driver"
            flavor        data
            legal_values  { 300 600 1200 2400 4800 9600 14400 19200 38400 
                            57600 115200 }
            default_value 38400
            description "
                This option specifies the default baud rate (speed) for the 
                eSCI port B."
        }

        cdl_option CYGNUM_IO_SERIAL_FREESCALE_ESCI_B_BUFSIZE {
            display       "Buffer size for the sSCI port A driver"
            flavor        data
            legal_values  0 to 8192
            default_value 128
            description   "
                This option specifies the size of the internal buffers used 
                for the eSCI port B."
        }
    
        cdl_option CYGNUM_IO_SERIAL_FREESCALE_ESCI_B_INT_PRIORITY {
            display      "eSCI prot B INTC priority"
            flavor       data
            legal_values 0 to 15
            default_value   7
            description "
                INTC has 16 interrupt levels: 0 (lowest) to 15 (highest).
            "
        }

    }

    cdl_component CYGPKG_IO_SERIAL_FREESCALE_ESCI_C {
        display       "eSCI port C driver"
        flavor        bool
        default_value 0
        description   "
            This option includes the serial device driver for the eSCI port C."

        cdl_option CYGDAT_IO_SERIAL_FREESCALE_ESCI_C_NAME {
            display       "Device name for eSCI port C"
            flavor        data
            default_value {"\"/dev/ser2\""}
            description   "
                This option specifies the device name for the eSCI port C."
        }

        cdl_option CYGNUM_IO_SERIAL_FREESCALE_ESCI_C_BAUD {
            display       "Baud rate for the eSCI serial port A driver"
            flavor        data
            legal_values  { 300 600 1200 2400 4800 9600 14400 19200 38400 
                            57600 115200 }
            default_value 38400
            description "
                This option specifies the default baud rate (speed) for the 
                eSCI port C."
        }

        cdl_option CYGNUM_IO_SERIAL_FREESCALE_ESCI_C_BUFSIZE {
            display       "Buffer size for the sSCI port A driver"
            flavor        data
            legal_values  0 to 8192
            default_value 128
            description   "
                This option specifies the size of the internal buffers used 
                for the eSCI port C."
        }
    
        cdl_option CYGNUM_IO_SERIAL_FREESCALE_ESCI_C_INT_PRIORITY {
            display      "eSCI prot B INTC priority"
            flavor       data
            legal_values 0 to 15
            default_value   6
            description "
                INTC has 16 interrupt levels: 0 (lowest) to 15 (highest).
            "
        }

    }

    cdl_component CYGPKG_IO_SERIAL_FREESCALE_ESCI_D {
        display       "eSCI port D driver"
        flavor        bool
        default_value 0
        description   "
            This option includes the serial device driver for the eSCI port D."

        cdl_option CYGDAT_IO_SERIAL_FREESCALE_ESCI_D_NAME {
            display       "Device name for eSCI port D"
            flavor        data
            default_value {"\"/dev/ser3\""}
            description   "
                This option specifies the device name for the eSCI port D."
        }

        cdl_option CYGNUM_IO_SERIAL_FREESCALE_ESCI_D_BAUD {
            display       "Baud rate for the eSCI serial port A driver"
            flavor        data
            legal_values  { 300 600 1200 2400 4800 9600 14400 19200 38400 
                            57600 115200 }
            default_value 38400
            description "
                This option specifies the default baud rate (speed) for the 
                eSCI port D."
        }

        cdl_option CYGNUM_IO_SERIAL_FREESCALE_ESCI_D_BUFSIZE {
            display       "Buffer size for the sSCI port A driver"
            flavor        data
            legal_values  0 to 8192
            default_value 128
            description   "
                This option specifies the size of the internal buffers used 
                for the eSCI port D."
        }
    
        cdl_option CYGNUM_IO_SERIAL_FREESCALE_ESCI_D_INT_PRIORITY {
            display      "eSCI prot B INTC priority"
            flavor       data
            legal_values 0 to 15
            default_value   6
            description "
                INTC has 16 interrupt levels: 0 (lowest) to 15 (highest).
            "
        }
    }


    cdl_component CYGPKG_IO_SERIAL_FREESCALE_ESCI_OPTIONS {
        display "Serial device driver build options"
        flavor  none
        description   "
            Package specific build options including control over
            compiler flags used only in building this package,
            and details of which tests are built."


        cdl_option CYGPKG_IO_SERIAL_FREESCALE_ESCI_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building these serial device drivers. These flags are
                used in addition to the set of global flags."
        }

        cdl_option CYGPKG_IO_SERIAL_FREESCALE_ESCI_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building these serial device drivers. These flags are
                removed from the set of global flags if present."
        }
    }
}

# EOF ser_freescale_esci.cdl
