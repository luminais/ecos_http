# ====================================================================
#
#      freebsd_net.cdl
#
#      Networking configuration data
#
# ====================================================================
# ####ECOSPDCOPYRIGHTBEGIN####                                    
# -------------------------------------------                     
# This file is part of eCos, the Embedded Configurable Operating System.
# Copyright (C) 2000, 2001, 2002 Free Software Foundation, Inc.   
#
# Permission is granted to use, copy, modify and redistribute this
# file.                                                           
#
# -------------------------------------------                     
# ####ECOSPDCOPYRIGHTEND####                                      
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      gthomas
# Original data:  gthomas
# Contributors:
# Date:           1999-11-29
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_NET_FREEBSD_STACK {
    display       "FreeBSD networking stack"
    parent        CYGPKG_NET
    doc           ref/tcpip-freebsd.html
    include_dir   .
    requires      CYGPKG_IO
    requires      CYGPKG_ISOINFRA
    requires      CYGINT_ISO_C_TIME_TYPES
    requires      CYGINT_ISO_STRERROR
    requires      CYGINT_ISO_ERRNO
    requires      CYGINT_ISO_ERRNO_CODES
    requires      CYGINT_ISO_MALLOC
    requires      CYGINT_ISO_STRING_BSD_FUNCS
    requires      CYGPKG_IO_FILEIO
    description   "Basic networking support, including TCP/IP."

    cdl_interface CYGINT_NET_IPSEC_BSD_CRYPTO {
        display   "Implementation of BSD CRYPTO functions"
        description "
          In order to avoid potential export problems of crypto
          functions, they are distributed in a separate package which
          must implement this interface"
    }

    implements    CYGPKG_NET_STACK
    implements    CYGPKG_NET_STACK_INET
    implements    CYGPKG_NET_STACK_INET6

    # Note: separating the stack implementation from the common support leads
    # to some rather incestious config file relationships.
    define_proc {
        puts $::cdl_system_header "/***** Networking stack proc output start *****/"
        puts $::cdl_header "#include <pkgconf/net.h>"
		#puts $::cdl_system_header "#define IPDIVERT 1"
	 	#puts $::cdl_system_header "#define IPFIREWALL 1"
	puts $::cdl_system_header "#define CYGDAT_NET_STACK_CFG <pkgconf/net_freebsd_stack.h>"
        puts $::cdl_system_header "/***** Networking stack proc output end *****/"
    }


    # Export our types to <sys/types.h>
    implements    CYGINT_ISO_BSDTYPES
    requires      { CYGBLD_ISO_BSDTYPES_HEADER == "<sys/bsdtypes.h>" }

    # These files are unique to eCos
    compile ecos/support.c \
        ecos/synch.c \
        ecos/timeout.c \
        ecos/init.cxx 
    compile -library=libextras.a sys/kern/sockio.c

    # These files were derived from FreeBSD and carry their copyright
    compile sys/net/if.c \
        sys/net/rtsock.c \
        sys/net/raw_cb.c \
        sys/net/raw_usrreq.c \
        sys/net/route.c \
        sys/net/radix.c \
        sys/net/if_ethersubr.c \
        sys/net/if_loop.c \
        sys/netinet/igmp.c \
        sys/netinet/raw_ip.c \
        sys/netinet/in.c  \
        sys/netinet/in_cksum.c \
        sys/netinet/in_pcb.c \
        sys/netinet/in_proto.c \
		sys/netinet/ip_gre.c \
        sys/netinet/in_rmx.c \
        sys/netinet/ip_encap.c \
        sys/netinet/ip_id.c \
        sys/netinet/ip_icmp.c \
        sys/netinet/ip_flow.c \
        sys/netinet/ip_input.c \
        sys/netinet/ip_output.c \
        sys/netinet/ip_mroute.c \
        sys/netinet/if_ether.c \
        sys/netinet/udp_usrreq.c \
        sys/netinet/tcp_input.c \
        sys/netinet/tcp_output.c \
        sys/netinet/tcp_debug.c \
        sys/netinet/tcp_usrreq.c \
        sys/netinet/tcp_timer.c \
        sys/netinet/tcp_subr.c \
        sys/kern/md5c.c \
        sys/kern/uipc_domain.c \
        sys/kern/uipc_socket.c \
        sys/kern/uipc_socket2.c \
        sys/kern/uipc_mbuf.c \
        sys/kern/uipc_mbuf2.c \
        sys/kern/uipc_accf.c \
        sys/kern/kern_subr.c

    cdl_component CYGPKG_NET_FREEBSD_PPPOE {
        display       "PPPOE support"
	active_if     CYGPKG_NET_INET 
	flavor	      bool
	define HAVE_PPPOE
	define HAVE_PPP_RTL
	default_value 0
	description    "
	    This option enables support for pppoe client processing."
	compile \
        	sys/net/pppoe.c \
	}

    cdl_component CYGPKG_NET_FREEBSD_L2TP {
        display       "L2TP support"
	active_if     CYGPKG_NET_INET 
	flavor	      bool
	define HAVE_L2TP
	define HAVE_PPP_RTL
	default_value 0
	description    "
	    This option enables support for l2tp client processing."
	compile \
        	sys/net/l2tp_avp_rtl.c \
        	sys/net/l2tp_ctrl_rtl.c \
        	sys/net/l2tp_rtl.c \
        	sys/net/l2tp_seq_rtl.c
	}

    cdl_component CYGPKG_NET_FREEBSD_DOUBLE_ALIAS {
        display       "double alias support"
        active_if     CYGPKG_NET_INET
        flavor        bool
        define CONFIG_RTL_SUPPORT_DOUBLE_ALIAS
        default_value 0
        description    "
            This option enables support for double alias."
        }

    cdl_component CYGPKG_NET_FREEBSD_PPTP {
        display       "PPTP support"
    active_if     CYGPKG_NET_INET
    flavor        bool
    define HAVE_PPTP
    default_value 0
    description    "
        This option enables support for pppt client processing."
    compile \
            sys/net/pptp/pptpd.c \
            sys/net/pptp/pptp_ctrl.c \
            sys/net/pptp/pptp_gre.c
    }

    cdl_component CYGPKG_NET_FREEBSD_NETGRAPH {
        display       "NETGRAPH support"
	active_if     CYGPKG_NET_INET 
	flavor	      bool
	define CYGPKG_NET_NETGRAPH
	default_value 0
	description    "
	    This option enables support for NEGGRAPH processing."
	compile \
		sys/netgraph/ng_base.c \
		sys/netgraph/ng_ether.c \
		sys/netgraph/ng_iface.c \
		sys/netgraph/ng_ksocket.c \
		sys/netgraph/ng_parse.c \
		sys/netgraph/ng_pppoe.c \
		sys/netgraph/ng_socket.c \
        	sys/kern/kern_module.c \
		sys/net/intrq.c
	}

    cdl_component CYGPKG_NET_FREEBSD_NETGRAPH_LIB {
        display       "NETGRAPH Library support"
        active_if     CYGPKG_NET_INET
        flavor        bool
        no_define
        default_value 0
        description    "
            This option enables support for NEGGRAPH library processing."
        compile \
                sys/libnetgraph/debug.c \
                sys/libnetgraph/msg.c \
                sys/libnetgraph/sock.c
        }
    cdl_component CYGPKG_NET_FREEBSD_INET {
        display       "INET support"
        active_if     CYGPKG_NET_INET
		flavor        bool
        no_define
        default_value 1
        description   "
            This option enables support for INET (IPv4) network processing."

		cdl_option CYGPKG_RTL_WANIP_SAME_WITH_GWIP_SUPPORT {
            display       "static or dhcp ip same with gateway support"
            default_value 0
            implements    CYGPKG_FREEBSD_RTL_WANIP_SAME_WITH_GWIP_SUPPORT
            flavor        bool

            description   "
                This option enables support for ip same with gw."
            # These files were derived from FreeBSD/KAME and carry their copyright
			define_proc {
		        puts $::cdl_system_header "#define CONFIG_RTL_WANIP_SAME_WITH_GWIP_SUPPORT 0"
    		}
        }
	
            cdl_option CYGPKG_RTL_DRV_DELIVER_INET {
            display       "driver deliver in inet"
            default_value 0
            implements    CYGPKG_FREEBSD_STACK_DRV_DELIVER_INET
            flavor        bool

            description   "
                This option enables support for drive deliver in inet thread."
            # These files were derived from FreeBSD/KAME and carry their copyright
                        define_proc {
                        puts $::cdl_system_header "#define CONFIG_RTL_DRV_DELIVER_INET 1"
                }
	}

		cdl_option CYGPKG_FAST_PATH {
            display       "fastpath support"
            default_value 0
            implements    CYGPKG_FREEBSD_STACK_FAST_PATH
            flavor        bool

            description   "
                This option enables support for fastpath."
            # These files were derived from FreeBSD/KAME and carry their copyright
			define_proc {
		        puts $::cdl_system_header "#define CONFIG_RTL_FREEBSD_FAST_PATH 0"
    		}
            compile \
                sys/netinet/fastpath/fastpath_core.S \
                sys/netinet/fastpath/fastpath_common.c \
				sys/netinet/fastpath/filter.S
        }

           cdl_option CYGPKG_FAST_PATH_PPPOE {
            display       "pppoe fastpath support"
            default_value 0
            implements    CYGPKG_FREEBSD_STACK_FAST_PATH
            flavor        bool

            description   "
                This option enables support for fastpath."
            # These files were derived from FreeBSD/KAME and carry their copyright
                        define_proc {
                        puts $::cdl_system_header "#define CONFIG_RTL_FAST_PPPOE 0"
                }
            compile \
                sys/netinet/fastpath/fast_pppoe_core.S 
        }	


			cdl_option CYGPKG_PPPOE_DIRECT_REPLY {
            display       "pppoe direct reply support"
            default_value 0
            implements    CYGPKG_FREEBSD_STACK_FAST_PATH
            flavor        bool
 
            description   "
                This option enables support for fastpath."
            # These files were derived from FreeBSD/KAME and carry their copyright
                        define_proc {
                        #puts $::cdl_system_header "#define CONFIG_RTL_PPPOE_DIRECT_REPLY 0"
                }
        	}

			cdl_option CYGPKG_FAST_PATH_L2TP {
            display       "L2TP fastpath support"
            default_value 0
            implements    CYGPKG_FREEBSD_STACK_FAST_PATH
            flavor        bool

            description   "
                This option enables support for fastpath."
            # These files were derived from FreeBSD/KAME and carry their copyright
                        define_proc {
                        puts $::cdl_system_header "#define FAST_L2TP 0"
                }
            compile \
                sys/netinet/fastpath/fast_l2tp_core.S
        	}
        
			cdl_option CYGPKG_FAST_PATH_PPTP {
			display       "PPTP fastpath support"
			default_value 0
			implements    CYGPKG_FREEBSD_STACK_FAST_PATH
            flavor        bool

			description   "
				This option enables support for fastpath."
			# These files were derived from FreeBSD/KAME and carry their copyright
						define_proc {
						puts $::cdl_system_header "#define FAST_PPTP 0"
			}
            compile \
                sys/netinet/fastpath/fast_pptp_core.S
        	}        
 	cdl_option CYGPKG_QOS_RATE_LIMIT_CHECK {
            display       "qos rate limit hook point"
            default_value 0
            implements    CYGPKG_FREEBSD_QOS_RATE_LIMIT_CHECK
            flavor        bool
            
            description   "
                This option enables for add hook point for qos rate limit."
            # These files were derived from FreeBSD/KAME and carry their copyright
                        define_proc {
                        puts $::cdl_system_header "#define CONFIG_RTL_QOS_RATE_LIMIT_CHECK 0"
                }       
        }       
    cdl_option CYGPKG_NAT_LOOPBACK {
            display       "nat loopback"
            default_value 0
            implements    CYGPKG_FREEBSD_NAT_LOOPBACK
            flavor        bool

            description   "
                This option enables for add nat loopback support."
            # These files were derived from FreeBSD/KAME and carry their copyright
                        define_proc {
                        puts $::cdl_system_header "#define CONFIG_RTL_NAT_LOOPBACK 0"
                }
        }
	cdl_option CYGPKG_NET_SNIPER {
            display       "bypass netsniper support"
            default_value 0
            implements    CYGPKG_FREEBSD_NET_SNIPER
            flavor        bool
 
            description   "
                This option enables support for bypass netsniper."
            # These files were derived from FreeBSD/KAME and carry their copyright
                        define_proc {
                        puts $::cdl_system_header "#define CONFIG_RTL_NETSNIPER_SUPPORT 0"
                }
            compile \
                sys/netinet/netsniper/rtl_netsniper.c
        }

	cdl_option CYGPKG_SPI_FIREWALL {
            display       "SPI(stateful packet inspection) firewall support"
            default_value 0
            implements    CYGPKG_FREEBSD_SPI_FIREWALL
            flavor        bool
 
            description   "
                This option enables support for SPI(stateful packet inspection) firewall."
            # These files were derived from FreeBSD/KAME and carry their copyright
                        define_proc {
                        puts $::cdl_system_header "#define CONFIG_RTL_SPI_FIREWALL_SUPPORT 0"
                }
            compile \
                sys/netinet/rtl_spi_firewall.c
        }

	cdl_option CYGPKG_FAST_PATH_SKB {
            display       "skb fastpath support"
            default_value 0
            implements    CYGPKG_FREEBSD_STACK_FAST_PATH_SKB
            flavor        bool
            description      "This option controls the skb fastpath" 
	    define_proc {
                        puts $::cdl_system_header "#define CONFIG_RTL_FREEBSD_FAST_PATH_SKB 0"
                }

	}
		cdl_option CYG_TCP_MAX_SOCKET_LIMITS {
		 display          "Maximum percentage of accept tcp socket"
        	 flavor           data
       		 default_value    2/3
       		 description      "This option controls the percentage of accept tcp socket
                          that if CONFIG_RTL_SORAPIDRECYCLE define"
               }

		 cdl_option CYGPKG_RTL_VLAN {
            display       "rtl vlan support"
            default_value 0
            implements    CYGPKG_FREEBSD_STACK_RTL_VLAN
            flavor        bool

            description   "
                This option enables support for rtl_vlan."
            # These files were derived from FreeBSD/KAME and carry their copyright
            define_proc {
                puts $::cdl_system_header "#define CONFIG_RTL_VLAN_SUPPORT 0"
            }
            compile \
                sys/netinet/rtl_vlan.c
		}		

		 cdl_option CYGPKG_RTL_BRIDGE_VLAN {
            display       "rtl bridge vlan support"
	    active_if     CYGPKG_RTL_VLAN 
            default_value 0
            implements    CYGPKG_FREEBSD_STACK_RTL_BRIDGE_VLAN
            flavor        bool

            description   "
                This option enables support for rtl bridge vlan."
            # These files were derived from FreeBSD/KAME and carry their copyright
            define_proc {
                puts $::cdl_system_header "#define CONFIG_RTL_BRIDGE_VLAN_SUPPORT 0"
            }
	    }

	    cdl_option CYGPKG_RTL_CONE_NAT {
            display       "rtl cone nat support"
	    	default_value 1
            implements    CYGPKG_FREEBSD_STACK_RTL_CONE_NAT
            flavor        bool

            description   "
                This option enables support for rtl_cone_nat."
            # These files were derived from FreeBSD/KAME and carry their copyright
            define_proc {
                puts $::cdl_system_header "#define CONFIG_RTL_CONE_NAT_SUPPORT 1"
            }
            compile \
                sys/netinet/libalias/alias_cone_nat.c
        }

		cdl_option CYGPKG_RTL_PORT_FWD {
           	display       "rtl port forwarding support"
        	default_value 1
            implements    CYGPKG_FREEBSD_STACK_RTL_PORT_FWD
            flavor        bool

            description   "
                This option enables support for rtl_port_fwd."
            # These files were derived from FreeBSD/KAME and carry their copyright
            define_proc {
                puts $::cdl_system_header "#define CONFIG_RTL_PORT_FORWARDING_SUPPORT 1"
            }
            compile \
                sys/netinet/libalias/alias_port_forwarding.c
        }

		cdl_option CYGPKG_RTL_TRIGGER_PORT {
            display       "rtl trigger port support"
            default_value 1
            implements    CYGPKG_FREEBSD_STACK_RTL_TRIGGER_PORT
            flavor        bool

            description   "
                This option enables support for rtl_trigger_port."
            # These files were derived from FreeBSD/KAME and carry their copyright
            define_proc {
                puts $::cdl_system_header "#define CONFIG_RTL_TRIGGER_PORT_SUPPORT 1"
            }
            compile \
                sys/netinet/libalias/alias_trigger_port.c
        }
	
		cdl_option CYGPKG_NET_FREEBSD_INET6 {
            display       "IPv6 support"
            active_if     CYGPKG_NET_INET6
            flavor        bool
            default_value 1
            description   "
                This option enables support for new IPv6."
            # These files were derived from FreeBSD and carry their copyright
            compile \
              sys/netinet6/dest6.c \
              sys/netinet6/frag6.c \
              sys/netinet6/icmp6.c \
              sys/netinet6/in6.c \
              sys/netinet6/in6_cksum.c \
              sys/netinet6/in6_ifattach.c \
              sys/netinet6/in6_pcb.c \
              sys/netinet6/in6_proto.c \
              sys/netinet6/in6_rmx.c \
              sys/netinet6/in6_src.c \
              sys/netinet6/ip6_forward.c \
              sys/netinet6/ip6_input.c \
              sys/netinet6/ip6_mroute.c \
              sys/netinet6/ip6_output.c \
              sys/netinet6/mld6.c \
              sys/netinet6/nd6.c \
              sys/netinet6/nd6_nbr.c \
              sys/netinet6/nd6_rtr.c \
              sys/netinet6/raw_ip6.c \
              sys/netinet6/route6.c \
              sys/netinet6/scope6.c \
              sys/netinet6/udp6_output.c \
              sys/netinet6/udp6_usrreq.c \

## Only if firewall enabled
##             sys/netinet6/ip6_fw.c \

        }

	cdl_component CYGPKG_NET_READYLOGO_PATCH {
       		display 	  "Patches for IPv6 ReadyLogo "
            active_if     CYGPKG_NET_INET6
			active_if 	  CYGPKG_NET_FREEBSD_INET6
			flavor 		  bool
            default_value 1
     		no_define
       		description "
              	This option controls IPv6 ReadyLogo patches support."

		cdl_option CYGPKG_NET_READYLOGO_CORE_PATCH {
            display       "IPv6 ReadyLogo Core patch"
            flavor        bool
            default_value 0
            description   "
                This option enables patches support for IPv6 ReadyLogo Core test."
        }
	}

	                cdl_option CYGPKG_FORWARD_FRAG_INET6 {
            display       "Forward ipv6 fragment support"
            flavor        bool
            default_value 0
            description   "
                This option enables patches support for Forward ipv6 fragment support."
        define_proc {
                puts $::cdl_system_header "#define CONFIG_FORWARD_IPV6_FRAG_SUPPORT 0"
        }
	}
        cdl_option CYGPKG_NET_FREEBSD_IPSEC {
            display       "IPSEC support"
            requires      CYGPKG_COMPRESS_ZLIB
            implements    CYGPKG_NET_STACK_IPSEC

            flavor        bool
            default_value CYGPKG_NET_IPSEC_BSD_CRYPTO

            description   "
                This option enables support for IPSEC."
            # These files were derived from FreeBSD/KAME and carry their copyright
            compile \
              sys/netkey/key.c \
              sys/netkey/key_debug.c \
              sys/netkey/keydb.c\
              sys/netkey/keysock.c \
              sys/netinet6/ipsec.c \
              sys/netinet6/ah_core.c \
              sys/netinet6/ah_input.c \
              sys/netinet6/ah_output.c \
              sys/netinet6/ipcomp_core.c \
              sys/netinet6/esp_core.c \
              sys/netinet6/esp_output.c \
              sys/netinet6/esp_input.c \
              sys/netinet6/esp_rijndael.c \
              sys/netinet6/esp_twofish.c \
              sys/netinet6/ipcomp_core.c \
              sys/netinet6/ipcomp_output.c \
              sys/netinet6/ipcomp_input.c \
              sys/netinet/ip_ecn.c
        }

	cdl_component CYGPKG_NET_BRIDGE {
         display "Built-in ethernet bridge code"
         default_value 0
         implements CYGINT_NET_BRIDGE_HANDLER
     	no_define
         description   "
             This option controls whether to include the built-in code for
             the Ethernet bridge."
     	compile sys/net/if_bridge.c 

         cdl_option CYGNUM_NET_BRIDGES {
             display "Number of Ethernet bridges"
             flavor  data
             default_value 1
             legal_values 1 to 999999
         }

         cdl_option CYGPKG_NET_BRIDGE_STP_CODE {
             display "Include code for Spanning Tree Protocol"
             default_value 0
             description "
                 This option controls whether to include the code for
                 the Spanning Tree Protocol on Ethernet bridge."
         }
    }
	
    cdl_interface CYGINT_NET_BRIDGE_HANDLER {
        display "Support for ethernet bridges in the IP stack"
        define NBRIDGE
            description "
              This interface controls whether calls to bridge code are made
              from the IP stack; these are needed if the built-in bridge code
              is used, but they can also be enabled in order to call different
              bridge code from an external component."
    }
	cdl_component CYGPKG_SAME_LAN_MAC {
       		display "Support eth0 and wlan0 with same mac address"
       		define CONFIG_SAME_LAN_MAC
       		description "
              	This option controls eth0 and wlan0 with same mac  support."
	}

    	cdl_component CYGPKG_NET_FIREWALL {
       		display "Support firewall"
       		define IPFIREWALL_FORWARD
		define_proc {
			puts $::cdl_system_header "#define IPFIREWALL 1"
       		}
		description "
              	This option controls firewall support."
			compile \
                        sys/netinet/ip_fw.c
	}

    	cdl_component CYGPKG_NET_IPV6FIREWALL {
       		display "Support ipv6 firewall"
       		define IPV6FIREWALL
       		define CONFIG_RTL_IPV6FIREWALL
       		description "
              	This option controls ipv6 firewall support."
			compile \
                        sys/netinet6/ip6_fw.c
	}
	cdl_component CYGPKG_NET_QOS {
       		display "Support QoS"
		active_if CYGPKG_NET_FIREWALL
		define DUMMYNET
       		description "
              	This option controls QoS support."
			compile \
			sys/netinet/ip_dummynet.c 
	}

	cdl_component CYGPKG_NET_NETBIOS {
       		display "Support NETBIOS"
			default_value 0
			define NETBIOS_SUPPORT
       		description "
              	This option controls NETBIOS support."
	}
	
	cdl_component CYGPKG_TIMER_HZ_1K {
            display       "Change HZ from 100 to 1000"
            define CYGPKG_TIMER_HZ_1K
            description   "
                This option change HZ to 1000"
    	}

	cdl_component CYGPKG_NET_IGMPPROXY_KERNEL_MODE {
    	display "igmp proxy kernel mode"
        default_value 0 
		define CONFIG_RTL_IGMP_PROXY_KERNEL_MODE
        define MROUTING    
        #description ""  
         }

 	cdl_component CYGPKG_NET_IGMPPROXY_USER_MODE {
    	display "igmp proxy user mode"
        default_value 0
        define CONFIG_RTL_IGMP_PROXY_USER_MODE
        define MROUTING
        #description ""
         }

	cdl_option CYGPKG_KLD_ENABLED {
			display "kld enable"
			default_value 0
			implements    CYGPKG_FREEBSD_STACK_KLD_ENABLED
            		flavor        bool
 
            		description   "
                	This option enables support for kld."
            		# These files were derived from FreeBSD/KAME and carry their copyright
                        define_proc {
                        puts $::cdl_system_header "#define KLD_ENABLED 0"
                }
	}

	cdl_component CYGPKG_NET_NAPT {
			display "Support napt"
			default_value 0
			define HAVE_NAPT
			define_proc {
				puts $::cdl_system_header "#define IPDIVERT 1"
			}
			description "
				This option controls napt support."
			compile \
				sys/netinet/ip_divert.c \
				sys/netinet/libalias/alias.c \
				sys/netinet/libalias/alias_cuseeme.c \
				sys/netinet/libalias/alias_db.c \
				sys/netinet/libalias/alias_nbt.c \
				sys/netinet/libalias/alias_proxy.c \
				sys/netinet/libalias/alias_util.c \
				sys/netinet/libalias/alias_irc.c \
				sys/netinet/libalias/alias_tftp.c \
				sys/netinet/libalias/alias_pptp_l2tp.c
	}

	cdl_component CYGPKG_NOT_NET_NATD {
                        display "Not support natd"
                        default_value 1
                        description "
                                This option controls not support natd."
        }	

	cdl_option CYGPKG_NET_KERNEL_NAPT {
            display       "Support kernel napt"
            active_if     CYGPKG_NET_NAPT
	    active_if	  CYGPKG_NOT_NET_NATD
            default_value 1
            description   "
                This option controls kernel napt support"
	
	    define_proc {
		puts $::cdl_system_header "#define CONFIG_RTL_NAPT_KERNEL_MODE_SUPPORT 1"
		#puts $::cdl_system_header "#define CONFIG_RTL_NAPT_TCP_GARBAGE_COLLECTION 1"
		#puts $::cdl_system_header "#define CONFIG_RTL_NAPT_GARBAGE_COLLECTION 1"
		}
            compile \
		sys/netinet/ip_napt.c
        }

	cdl_component CYGPKG_NET_NAT_ALG {
			display "Support nat alg"
            		active_if CYGPKG_NET_NAPT
			default_value 0
			define HAVE_NAT_ALG
			description "
				This option controls nat alg support."
	}
        cdl_option CYGPKG_NET_NAT_ALG_FTP {
            display       "Support ftp alg"
            active_if	  CYGPKG_NET_NAPT
            active_if	  CYGPKG_NET_NAT_ALG
            default_value 1
	    define HAVE_NAT_ALG_FTP
            description   "
                This option controls ftp alg support"

            compile \
              sys/netinet/libalias/alias_ftp.c 
        } 
        cdl_option CYGPKG_NET_NAT_ALG_RTSP {
            display       "Support rtsp alg"
            active_if	  CYGPKG_NET_NAPT
            active_if	  CYGPKG_NET_NAT_ALG
            default_value 1
	    define HAVE_NAT_ALG_RTSP
            description   "
                This option controls rtsp alg support"

            compile \
              sys/netinet/libalias/alias_smedia.c
        } 
        cdl_option CYGPKG_NET_NAT_ALG_SIP {
            display       "Support sip alg"
            active_if	  CYGPKG_NET_NAPT
            active_if	  CYGPKG_NET_NAT_ALG
            default_value 1
	    define HAVE_NAT_ALG_SIP
            description   "
                This option controls sip alg support"

            compile \
              sys/netinet/libalias/alias_sip.c
        } 
        cdl_option CYGPKG_NET_NAT_ALG_PPTP {
            display       "Support pptp alg"
            active_if	  CYGPKG_NET_NAPT
            active_if	  CYGPKG_NET_NAT_ALG
            default_value 1
	    define HAVE_NAT_ALG_PPTP
            description   "
                This option controls pptp alg support"
        } 
        cdl_option CYGPKG_NET_NAT_ALG_L2TP {
            display       "Support l2tp alg"
            active_if	  CYGPKG_NET_NAPT
            active_if	  CYGPKG_NET_NAT_ALG
            default_value 1
	    define HAVE_NAT_ALG_L2TP
            description   "
                This option controls l2tp alg support"
        } 
        cdl_option CYGPKG_NET_NAT_ALG_TFTP {
            display       "Support tftp alg"
            active_if	  CYGPKG_NET_NAPT
            active_if	  CYGPKG_NET_NAT_ALG
            default_value 1
	    define HAVE_NAT_ALG_TFTP
            description   "
                This option controls tftp alg support"

            compile \
              sys/netinet/libalias/alias_tftp.c
        } 
	cdl_option CYGPKG_NET_NAT_ALG_H323 {
            display       "Support h323 alg"
            active_if     CYGPKG_NET_NAPT
            active_if     CYGPKG_NET_NAT_ALG
            default_value 0
            define HAVE_NAT_ALG_H323
            description   "
                This option controls h323 alg support"
 
            compile \
	      sys/netinet/libalias/alias_h323_asn1.c \
	      sys/netinet/libalias/alias_h323_main.c
        }

    cdl_option CYGPKG_NET_FREEBSD_IPSEC6 {
            display       "IPSEC support for IPv6"
            active_if     CYGPKG_NET_INET6
            active_if     CYGPKG_NET_FREEBSD_IPSEC

            flavor        bool
            default_value 1
            description   "
                This option enables support for IPSEC with IPv6"
            compile \
              sys/netinet6/in6_gif.c

        }
        cdl_option CYGPKG_NET_FREEBSD_SYSCTL {
            display       "sysctl support"
            flavor        bool
            default_value 1
            description   "
                This option enables support for the system call sysctl used
            to configure options/variables in the stack and retrieve statistics. "
            # This file was derived from FreeBSD and carries that copyright
            compile \
              sys/kern/kern_sysctl.c
        } 
        cdl_option CYGPKG_NET_RANDOM_PORTS {
            display       "Random source ports"
            flavor        bool
            default_value 0
            description   "
                This option enables support for random source ports when the source
            port is not specified.  This option is useful when connecting
            through firewalls."
        }                 
    }

    cdl_option CYGPKG_NET_NGIF {
        display "Number of GIF things"
        flavor  data
        default_value 0
        description   "
            This option controls the number of active GIF things."
        define NGIF
    }

    cdl_option CYGPKG_NET_NLOOP {
        display "Number of loopback interfaces"
        flavor  data
        default_value 1
        description   "
            This option controls the number of loopback, i.e. local, interfaces.
            There is seldom need for this value to be anything other than one."
        define NLOOP
    }

    cdl_option CYGPKG_NET_FREEBSD_LOGGING {
        display       "Error and warning log control"
        flavor        booldata
        default_value 0xC08F
        description   "
            This option controls the type and amount of information
            printed by the networking code.  Different logging 
            facilities may be enabled by bitwise or-ing:
              LOG_ERR     0x0001 - error conditions
              LOG_WARNING 0x0002 - interesting, but not errors
              LOG_NOTICE  0x0004 - things to look out for
              LOG_INFO    0x0008 - generic comments
              LOG_DEBUG   0x0010 - for finding obscure problems
              LOG_MDEBUG  0x0020 - additional information about memory allocations
              LOG_IOCTL   0x0040 - information about ioctl calls
              LOG_INIT    0x0080 - information as system initializes
              LOG_ADDR    0x0100 - information about IPv6 addresses
              LOG_FAIL    0x0200 - why packets (IPv6) are ignored, etc.
              LOG_EMERG   0x4000 - emergency conditions
              LOG_CRIT    0x8000 - critical error
            "
    }

    cdl_option CYGPKG_NET_FORCE_SERIAL_CONSOLE {
        display "Force use of serial console during initialization"
        flavor  bool
        default_value 0
        description   "
            Trying to print initialization messages can fail if the
            console channel is a network connection (via RedBoot).
            Use of this option forces the stack to use a serial
            port during this phase for safety.  It can be used 
            if the network drivers are unstable at this point."
    }

    cdl_option CYGPKG_NET_MEM_USAGE {
        display "Memory designated for networking buffers."
        flavor  data
        default_value (256*1024)+(CYGPKG_NET_MAXSOCKETS*1024)
        description   "
            This option controls the amount of memory pre-allocated
        for buffers used by the networking code.  The number is an
        upper limit, with at least enough space to get the stack
        initialized. Tip: setting a breakpoint at cyg_memalloc_alloc_fail() 
	is an especially useful tool in establishing when there is too 
        little memory for an application. "
    }

    cdl_option CYGPKG_NET_MEMPOOL_SIZE {
        display "Memory designated for network dynamically allocated memory"
        flavor  data
        default_value CYGPKG_NET_MEM_USAGE/4
        description   "
            Controls the amount of memory in the pool used for dynamically
            allocated memory. This does not include mbufs or clusters."
    }

    cdl_option CYGPKG_NET_MBUFS_SIZE {
        display "MBUFs memory size"
        flavor  data
        default_value CYGPKG_NET_MEM_USAGE/4
        description   "
            Size of MBUFs pool."
    }

    cdl_option CYGPKG_NET_CLUSTERS_SIZE {
        display "Clusters size"
        flavor  data
        default_value CYGPKG_NET_MEM_USAGE/2
        description   "
            Clusters size."
    }

    cdl_option CYGPKG_NET_MAXSOCKETS {
        display "Max number of open sockets"
        flavor  data
        default_value CYGNUM_FILEIO_NFILE
        description   "
            This option controls the amount of memory pre-allocated
        for socket buffers used by the networking code."
    }

    cdl_option CYGPKG_NET_NUM_WAKEUP_EVENTS {
        display "Number of supported pending network events"
        flavor  data
        default_value 8
        description   "
            This option controls the number of pending network events
        used by the networking code."
    }

    cdl_component CYGPKG_NET_THREAD {
        display        "Background network processing thread options"
        flavor        none
        no_define

     cdl_option CYGPKG_NET_THREAD_PRIORITY {
            display "Priority level for background network processing"
            flavor  data
            default_value 7
            description   "
                This option allows the thread priority level used by the
            networking stack to be adjusted by the user.  It should be set
            high enough that sufficient CPU resources are available to
            process network data, but may be adjusted so that application
            threads can have precedence over network processing."
        }

        cdl_option CYGNUM_NET_THREAD_STACKSIZE {
            display "Stack size for backgound network processing"
            flavor  data
            default_value { (CYGPKG_NET_INET6 ? 
                             "CYGNUM_HAL_STACK_SIZE_TYPICAL+2048" :
                             "CYGNUM_HAL_STACK_SIZE_TYPICAL") }
            description   "
                This option allows the thread stack allocated for the
            networking stack to be adjusted by the user. "
        }
    }

    cdl_component CYGPKG_NET_FAST_THREAD {
        display       "Fast network processing thread options"
        flavor        none
        no_define

        cdl_option CYGPKG_NET_FAST_THREAD_PRIORITY {
            display       "Priority level for fast network processing"
            flavor        data
            default_value CYGPKG_NET_THREAD_PRIORITY - 1
            description   "
                This option sets the thread priority level used by the fast
            network thread.  The fast network thread runs often but briefly, to
            service network device interrupts and network timeout events.  This
            thread should have higher priority than the background network
            thread.  It is reasonable to set this thread's priority higher than
            application threads for best network throughput, or to set it lower
            than application threads for best latency for those application
            threads themselves, potentially at a cost to network throughput."
        }

        cdl_option CYGNUM_NET_FAST_THREAD_STACKSIZE {
            display       "Stack size for fast network processing"
            flavor        data
            default_value { "CYGNUM_HAL_STACK_SIZE_TYPICAL" }
            description   "
                This option allows the thread stack allocated for the
            fast networking stack to be adjusted by the user. "
        }
    }

    cdl_component CYGPKG_NET_FAST_THREAD_TICKLE_DEVS {
        display "Fast network processing thread 'tickles' drivers"
        default_value 1
        description "
            If this is enabled, the fast network thread will tickle the
            device(s) periodically, to unblock them when the hardware has
            become wedged due to a lost interrupt or other hardware
            race-condition type problem.
            This is not necessary if a networked app is running which sends
            packets itself often - or
            uses TCP, or any similar protocol which exchanges keep-alive
            packets periodically and often enough.
            Trying to send a packet passes control into the driver; this is
            sufficient to detect and unblock jammed hardware."

        cdl_option CYGNUM_NET_FAST_THREAD_TICKLE_DEVS_DELAY {
            display "Delay in kernel clocks of tickle loop"
            flavor data
            default_value 50
            description "
                The default is 50, which will usually mean a delay between
                tests for 'stuck' devices of 500mS, that is half a second.
	        The overhead only applies if no network activity occurred,
	        so it may be acceptable to make this value very small,
                where high CPU load does not matter during network idle
                periods, or very large if your application tries often to
                send packets itself."
        }
    }

    cdl_component CYGPKG_NET_FREEBSD_STACK_OPTIONS {
        display "Networking support build options"
        flavor  none
        no_define

        cdl_option CYGOPT_NET_FREEBSD_STACK_ACCEPT_UNICAST {
            display "Accept unicast packets on INADDR_ANY interfaces"
            flavor  bool
            no_define
            define        BOOTP_COMPAT
            default_value 0
            description   "This option enables passing of unicast
                IP packets to the application, when the interface
                IP address is configured as INADDR_ANY (0.0.0.0).
                This option is useful for some applications that
                need to receive unicast IP packets when the interface
                address is unknown.  Such an application is bootp."
        }

        cdl_option CYGPKG_NET_FREEBSD_STACK_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { ( CYGPKG_NET_INET6? "-D_KERNEL -DGATEWAY6" : "-D_KERNEL" ) }
            description   "
                This option modifies the set of compiler flags for
                building the networking package.
                These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_NET_FREEBSD_STACK_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the networking package. These flags are removed from
                the set of global flags if present."
        }
    }
    cdl_option CYGPKG_NET_FREEBSD_STACK_TESTS {
        display       "FreeBSD network stack tests"
        flavor        data
        no_define
        calculated { CYGPKG_NET_FREEBSD_SYSCTL ? "tests/sysctl1" : "" }
        description  "
            These are test specifically for the FreeBSD stack. These test features
            which only the FreeBSD stack has"
    }
    cdl_option CYGPKG_NET_FREEBSD_MBUF_SHRINK {
        display       "FreeBSD network mbuf usage reduce"
        flavor        data
        define RTL_SMALL_MBUF
        description  "
            These are specifically for the FreeBSD stack. These test features
            which only the FreeBSD stack has"
    }

   cdl_option CYGPKG_NET_FREEBSD_GET_MEMINFO {
        display         "Display Miscpool and cluster size"
        flavor          bool
        default_value   0
        description     "
                This gives the mem chain upgrade support when update firemare."
    }
}
