# ====================================================================
#
#      flash_edb7xxx.cdl
#
#      FLASH memory - Hardware support on Cirrus Logic EDB7xxx
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      gthomas
# Original data:  gthomas
# Contributors:
# Date:           2000-07-26
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_FLASH_EDB7XXX {
    display       "FLASH support for Cirrus Logic EP7xxx based boards"
    description   "FLASH memory device support for Cirrus Logic EP7xxx based 
                   development boards"

    parent        CYGPKG_IO_FLASH
    active_if	  CYGPKG_IO_FLASH
    requires	  CYGPKG_HAL_ARM_EDB7XXX
    include_dir   cyg/io

    cdl_component CYGPKG_DEVS_FLASH_EP72XX {
        display       "Cirrus Logic EP72xx based boards"
        description    "FLASH memory device support for EP72xx based boards
                        specifically"
        active_if     { CYGHWR_HAL_ARM_EDB7XXX_BOARD_VARIANT != "EDB7312" }
        calculated    1
        no_define
        implements    CYGHWR_IO_FLASH_DEVICE
        implements    CYGHWR_IO_FLASH_DEVICE_LEGACY
    
        compile       edb7xxx_flash.c flash_query.c flash_program_buf.c flash_erase_block.c
    
    }
    cdl_component CYGPKG_DEVS_FLASH_STRATA_EDB7XXX {
        display       "Cirrus Logic EDB7xxx StrataFLASH memory support"
        description   "FLASH memory device support for Cirrus Logic EP73xx"
    
        # Note: currently only available on 7312 boards
        active_if     { CYGHWR_HAL_ARM_EDB7XXX_BOARD_VARIANT == "EDB7312" }
        requires      CYGPKG_DEVS_FLASH_STRATA
        calculated    1
        no_define    
    
        implements    CYGHWR_IO_FLASH_BLOCK_LOCKING
    
        # Arguably this should do in the generic package
        # but then there is a logic loop so you can never enable it.
        cdl_interface CYGINT_DEVS_FLASH_STRATA_REQUIRED {
            display   "Generic StrataFLASH driver required"
        }
    
        implements    CYGINT_DEVS_FLASH_STRATA_REQUIRED
    
        define_proc {
            puts $::cdl_system_header "/***** strataflash driver proc output start *****/"
            puts $::cdl_system_header "#define CYGDAT_DEVS_FLASH_STRATA_INL <cyg/io/edb7xxx_strataflash.inl>"
            puts $::cdl_system_header "#define CYGDAT_DEVS_FLASH_STRATA_CFG <pkgconf/devs_flash_edb7xxx.h>"
            puts $::cdl_system_header "/*****  strataflash driver proc output end  *****/"
        }
    }
}
