# ====================================================================
#
#      hal_powerpc_quicc.cdl
#
#      PowerPC/QUICC HAL package configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002, 2003 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Original data:  hmt
# Contributors:
# Date:           1999-11-02
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_QUICC {
    display  "Motorola MPC8xx PowerQUICC support"
    parent        CYGPKG_HAL_POWERPC
    define_header hal_powerpc_quicc.h
    include_dir   cyg/hal/quicc
    description   "
           The QUICC package provides some of the support needed
           to run eCos on a Motorola MPC8xx (MBX) board, using the QUICC
           feature of the MPC860 and MPC821 CPUs.
           Currently only serial IO via SMC1/2 and SCC1 is provided by
           this package."

    define_proc {
        puts $::cdl_system_header "#define CYGBLD_HAL_VARIANT_H  <pkgconf/hal_powerpc_quicc.h>"
    }

    cdl_interface CYGNUM_HAL_QUICC_SMC1 {
        display    "SMC1 is available for serial I/O"
        description "
          This interface indicates that SMC1 can be outfitted as
          a serial device."
    }

    cdl_interface CYGNUM_HAL_QUICC_SMC2 {
        display    "SMC2 is available for serial I/O"
        description "
          This interface indicates that SMC2 can be outfitted as
          a serial device."
    }

    cdl_interface CYGNUM_HAL_QUICC_SCC1 {
        display    "SCC1 is available for serial I/O"
        description "
          Most MPC8xx chipsets use SCC1 to drive the ethernet controller.
        On some newer (e.g. 860T) chips, SCC1 can be used for general
        serial since there is a separate ethernet machine."
    }

    cdl_interface CYGNUM_HAL_QUICC_SCC2 {
        display    "SCC2 is available for serial I/O"
        description "
          Port SCC2 is available for serial I/O"
    }

    cdl_interface CYGNUM_HAL_QUICC_SCC3 {
        display    "SCC3 is available for serial I/O"
        description "
          Port SCC3 is available for serial I/O"
    }

    cdl_interface CYGNUM_HAL_QUICC_SCC4 {
        display    "SCC4 is available for serial I/O"
        description "
          Port SCC4 is available for serial I/O"
    }

    compile       quicc_smc1.c cpm.c

   cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS {
       display      "Number of communication channels on the board"
       flavor       data
       calculated   CYGNUM_HAL_QUICC_SMC1+CYGNUM_HAL_QUICC_SMC2+CYGNUM_HAL_QUICC_SCC1+CYGNUM_HAL_QUICC_SCC2+CYGNUM_HAL_QUICC_SCC3+CYGNUM_HAL_QUICC_SCC4
   }

   cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL {
       display          "Debug serial port"
       active_if        CYGPRI_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_CONFIGURABLE
       flavor data
       legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
       default_value    0
       description      "
           This option chooses which port will be used to connect to a host
           via the GDB remote protocol."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL {
        display          "Diagnostic serial port"
        active_if        CYGPRI_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_CONFIGURABLE
        flavor data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        default_value    0
        description      "
           This option chooses which port will be used for diagnostic output."
    }

    # This option is only used when USE_ROM_MONITOR is enabled - but
    # it cannot be a sub-option to that option, since the code uses the
    # definition in a preprocessor comparison.
    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_ROM_DEBUG_CHANNEL {
        display          "Debug serial port used by ROM monitor"
        flavor data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        default_value    0
        description      "
            If a platform has multiple serial ports, then this
            option tells the code which port is in use by the ROM
            monitor. It should only be necessary to change this
            option if a non-standard configurated eCos GDB stub is
            used."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_BAUD {
        display       "Baud rate for the HAL diagnostic port"
        flavor        data
        legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                      4800 7200 9600 14400 19200 38400 57600 115200 230400
        }
        default_value 38400
        description   "
            This option specifies the default baud rate (speed) for the 
            HAL diagnostic port."
    }

}
