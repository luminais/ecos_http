# ====================================================================
#
#      linux.cdl
#
#      Linux compatibility layer data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002, 2003 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      dwmw2
# Contributors:   tkoeller
# Date:           2003-01-08
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_LINUX_COMPAT {
    display       "Linux compatibility layer"
    include_dir   ""
    description   "
	eCos supports a basic Linux compatibility Layer providing various
        functions, equivalents or stubs expected by Linux kernel code, for
        assistance in porting drivers and file system code from Linux.
        Note this does not provide Linux compatibility to applications."

    compile      rbtree.c

    cdl_option CYGNUM_LINUX_COMPAT_PAGE_SIZE_EXPONENT {
        display         "Define page size"
        flavor          data
        legal_values    10 to 16
        default_value   12
        no_define
        define          PAGE_SHIFT
        description     "
            Define the page size. The value entered here is used as an
            exponent X in the expression 2^^X to ensure that the page
            size is always an integer power of two."  
     } 
}

# EOF linux.cdl
