# ====================================================================
#
#      ser_i386_pc.cdl
#
#      eCos serial PC configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jlarmour, nickg, gthomas, pjo
# Original data:  
# Contributors:   jskov
# Date:           2001-06-08
#
#####DESCRIPTIONEND####
#
# ====================================================================


cdl_package CYGPKG_IO_SERIAL_I386_PC {
    display       "PC serial device drivers"

    parent        CYGPKG_IO_SERIAL_DEVICES
    active_if     CYGPKG_IO_SERIAL
    active_if     CYGPKG_HAL_I386_PCMB

    requires      CYGPKG_ERROR
    include_dir   cyg/io
    description   "
           This option enables the serial device drivers for the
           PC."

    # FIXME: This really belongs in the GENERIC_16X5X package
    cdl_interface CYGINT_IO_SERIAL_GENERIC_16X5X_REQUIRED {
        display   "Generic 16x5x serial driver required"
    }

    define_proc {
        puts $::cdl_system_header "/***** serial driver proc output start *****/"
        puts $::cdl_system_header "#define CYGDAT_IO_SERIAL_GENERIC_16X5X_INL <cyg/io/i386_pc_ser.inl>"
        puts $::cdl_system_header "#define CYGDAT_IO_SERIAL_GENERIC_16X5X_CFG <pkgconf/io_serial_i386_pc.h>"
        puts $::cdl_system_header "/*****  serial driver proc output end  *****/"
    }

cdl_component CYGPKG_IO_SERIAL_I386_PC_SERIAL0 {
    display       "PC serial port 0 driver"
    flavor        bool
    default_value 1
    description   "
        This option includes the serial device driver for port 0 on the 
        PC."

    implements    CYGINT_IO_SERIAL_GENERIC_16X5X_REQUIRED
    implements    CYGINT_IO_SERIAL_FLOW_CONTROL_HW
    implements    CYGINT_IO_SERIAL_LINE_STATUS_HW

    cdl_option CYGDAT_IO_SERIAL_I386_PC_SERIAL0_NAME {
        display       "Device name for PC serial port 0"
        flavor        data
        default_value {"\"/dev/ser0\""}
        description   "
            This option specifies the device name port 0 on the PC."
    }

    cdl_option CYGNUM_IO_SERIAL_I386_PC_SERIAL0_BAUD {
        display       "Baud rate for the PC serial port 0 driver"
        flavor        data
        legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                      4800 7200 9600 14400 19200 38400 57600 115200 230400
        }
        default_value 38400
        description   "
            This option specifies the default baud rate (speed) for the
            PC port 0."
    }

    cdl_option CYGNUM_IO_SERIAL_I386_PC_SERIAL0_BUFSIZE {
        display       "Buffer size for the PC serial port 0 driver"
        flavor        data
        legal_values  0 to 8192
        default_value 128
        description   "
            This option specifies the size of the internal buffers used
            for the PC port 0."
    }

    cdl_option CYGNUM_IO_SERIAL_I386_PC_SERIAL0_IOBASE {
	display "I/O base address for the i386-PC serial port 0"
	flavor    data
	legal_values 0 to 0xFF8
	default_value 0x3F8
	description "
	This option specifies the I/O address of the 8250 or 16550 for serial port 0."
    }

    cdl_option CYGNUM_IO_SERIAL_I386_PC_SERIAL0_IRQ {
	display "IRQ for the i386-PC serial port 0"
	flavor    data
	legal_values 0 to 15
	default_value 4
	description "
	This option specifies the IRQ of the 8250 or 16550 for serial port 0."
   }

    cdl_option CYGNUM_IO_SERIAL_I386_PC_SERIAL0_INT {
	display "INT for the i386-PC serial port 0"
	flavor    data
	legal_values 32 to 47
	default_value { CYGNUM_IO_SERIAL_I386_PC_SERIAL0_IRQ + 32 }
	description "
	This option specifies the interrupt vector of the 8250 or 16550 for serial port 0."
   }
}

cdl_component CYGPKG_IO_SERIAL_I386_PC_SERIAL1 {
    display       "PC serial port 1 driver"
    flavor        bool
    default_value 1
    description   "
        This option includes the serial device driver for port 1 on
        the PC."

    implements    CYGINT_IO_SERIAL_GENERIC_16X5X_REQUIRED
    implements    CYGINT_IO_SERIAL_FLOW_CONTROL_HW
    implements    CYGINT_IO_SERIAL_LINE_STATUS_HW

    cdl_option CYGDAT_IO_SERIAL_I386_PC_SERIAL1_NAME {
        display       "Device name for PC serial port 1"
        flavor        data
        default_value {"\"/dev/ser1\""}
        description   "
            This option specifies the device name port 1 on the PC."
    }

    cdl_option CYGNUM_IO_SERIAL_I386_PC_SERIAL1_BAUD {
        display       "Baud rate for the PC serial port 1 driver"
        flavor        data
        legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                      4800 7200 9600 14400 19200 38400 57600 115200 230400
        }
        default_value 38400
        description   "
            This option specifies the default baud rate (speed) for the
	    PC port 1."
    }

    cdl_option CYGNUM_IO_SERIAL_I386_PC_SERIAL1_BUFSIZE {
        display       "Buffer size for the PC serial port 1 driver"
        flavor        data
        legal_values  0 to 8192
        default_value 128
        description   "
            This option specifies the size of the internal buffers used
	    for the PC port 1."
    }

    cdl_option CYGNUM_IO_SERIAL_I386_PC_SERIAL1_IOBASE {
	display "I/O base address for the i386-PC serial port 1"
	flavor    data
	legal_values 0 to 0xFF8
	default_value 0x2F8
	description "
	This option specifies the I/O address of the 8250 or 16550 for serial port 1."
    }

    cdl_option CYGNUM_IO_SERIAL_I386_PC_SERIAL1_IRQ {
	display "IRQ for the i386-PC serial port 1"
	flavor    data
	legal_values 0 to 15
	default_value 3
	description "
	This option specifies the IRQ of the 8250 or 16550 for serial port 1."
   }

    cdl_option CYGNUM_IO_SERIAL_I386_PC_SERIAL1_INT {
	display "INT for the i386-PC serial port 1"
	flavor    data
	legal_values 32 to 47
	default_value { CYGNUM_IO_SERIAL_I386_PC_SERIAL1_IRQ + 32 }
	description "
	This option specifies the interrupt vector of the 8250 or 16550 for serial port 1."
   }
}

    cdl_component CYGPKG_IO_SERIAL_I386_PC_OPTIONS {
        display "Serial device driver build options"
        flavor  none
        description   "
	    Package specific build options including control over
	    compiler flags used only in building this package,
	    and details of which tests are built."


        cdl_option CYGPKG_IO_SERIAL_I386_PC_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building these serial device drivers. These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_IO_SERIAL_I386_PC_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building these serial device drivers. These flags are removed from
                the set of global flags if present."
        }
    }

    cdl_component CYGPKG_IO_SERIAL_I386_PC_TESTING {
        display    "Testing parameters"
        flavor     bool
        calculated 1
        active_if  CYGPKG_IO_SERIAL_I386_PC_SERIAL0

        cdl_option CYGPRI_SER_TEST_SER_DEV {
            display       "Serial device used for testing"
            flavor        data
            default_value { CYGDAT_IO_SERIAL_I386_PC_SERIAL0_NAME }
        }

        define_proc {
            puts $::cdl_header "#define CYGPRI_SER_TEST_CRASH_ID \"i386pc\""
            puts $::cdl_header "#define CYGPRI_SER_TEST_TTY_DEV  \"/dev/tty0\""
        }
    }
}

# EOF ser_i386_pc.cdl
