# ====================================================================
#
#      edosk2674_eth_drivers.cdl
#
#      Ethernet drivers - support for LAN91CXX ethernet controller
#      on the EDOSK-2674 board.
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      yoshinori sato
# Contributors:   yoshinori sato
# Date:           2003-02-26
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_ETH_H8300_EDOSK2674 {

    display       "EDOSK-2674 SMC91C96 ethernet driver"

    parent        CYGPKG_IO_ETH_DRIVERS
    active_if	  CYGPKG_IO_ETH_DRIVERS
    active_if	  CYGPKG_HAL_H8300_H8S_EDOSK2674

    implements    CYGHWR_NET_DRIVERS
    implements    CYGHWR_NET_DRIVER_ETH0
    implements    CYGINT_DEVS_ETH_SMSC_LAN91CXX_REQUIRED
    implements    CYGSEM_DEVS_ETH_SMSC_LAN91CXX_8_BIT

    description   "Ethernet driver for EDOSK-2674 boards."

    include_dir   cyg/io

    define_proc {
        puts $::cdl_system_header "/***** ethernet driver proc output start *****/"
        puts $::cdl_system_header "#define CYGDAT_DEVS_ETH_SMSC_LAN91CXX_INL <cyg/io/devs_eth_edosk2674.inl>"
        puts $::cdl_system_header "#define CYGDAT_DEVS_ETH_SMSC_LAN91CXX_CFG <pkgconf/devs_eth_h8300_edosk2674.h>"
        puts $::cdl_system_header "/*****  ethernet driver proc output end  *****/"
    }
    
    # Arguably this should do in the generic package
    # but then there is a logic loop so you can never enable it.

    cdl_interface CYGINT_DEVS_ETH_SMSC_LAN91CXX_REQUIRED {
        display   "SMSC LAN91CXX driver required"
    }

    cdl_option CYGDAT_DEVS_ETH_H8300_EDOSK2674_NAME {
        display       "Device name for the ethernet driver"
        flavor        data
        default_value {"\"eth0\""}
        description   "
            This option sets the name of the ethernet device for the
            ethernet port."
    }

    cdl_option CYGDAT_DEVS_ETH_H8300_EDOSK2674_ESA {
        display       "The ethernet station address (MAC)"
        flavor        data
        default_value {"{0x12, 0x13, 0x14, 0x15, 0x16, 0x17}"}
        description   "A static ethernet station address. 
            Caution: Booting two systems with the same MAC on the same
            network, will cause severe conflicts."
        active_if     !CYGSEM_DEVS_ETH_ARM_FLEXANET_REDBOOT_ESA
    }

    cdl_option CYGSEM_DEVS_ETH_H8300_EDOSK2674_ETH0_SET_ESA {
        display "Use the RedBoot ESA (MAC address)"
        default_value 0
        flavor        bool
        description   "
            Use the ESA that is stored as a RedBoot variable instead of
            a static ESA." 
    }

}

# EOF flexanet_eth_drivers.cdl
