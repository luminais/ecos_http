# ====================================================================
#
#      ser_arm_cerfpda.cdl
#
#      eCos serial CERFPDA configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Original data:  gthomas
# Contributors:
# Date:           1999-07-07
#
#####DESCRIPTIONEND####
#
# ====================================================================


cdl_package CYGPKG_IO_SERIAL_ARM_CERFPDA {
    display       "Cerfpda 16x5x serial device driver"

    parent        CYGPKG_IO_SERIAL_DEVICES
    active_if     CYGPKG_IO_SERIAL
    active_if     CYGPKG_HAL_ARM_SA11X0_CERFPDA

    requires      CYGPKG_ERROR
    include_dir   cyg/io

    description   "
           This option enables the serial 16x5x device drivers for the
           Cerfpda."

    # FIXME: This really belongs in the GENERIC_16X5X package
    cdl_interface CYGINT_IO_SERIAL_GENERIC_16X5X_REQUIRED {
        display   "Generic 16x5x serial driver required"
    }
    define_proc {
        puts $::cdl_header "#define CYGPRI_IO_SERIAL_GENERIC_16X5X_STEP 4"
    }


    define_proc {
        puts $::cdl_system_header "/***** serial driver proc output start *****/"
        puts $::cdl_system_header "#define CYGDAT_IO_SERIAL_GENERIC_16X5X_INL <cyg/io/arm_sa11x0_cerfpda_ser.inl>"
        puts $::cdl_system_header "#define CYGDAT_IO_SERIAL_GENERIC_16X5X_CFG <pkgconf/io_serial_arm_cerfpda.h>"
        puts $::cdl_system_header "/*****  serial driver proc output end  *****/"
    }


    cdl_component CYGPKG_IO_SERIAL_ARM_CERFPDA_SERIAL1 {
        display       "Cerfpda serial port 1 driver"
        flavor        bool
        default_value 1

        implements CYGINT_IO_SERIAL_GENERIC_16X5X_REQUIRED
        implements CYGINT_IO_SERIAL_FLOW_CONTROL_HW
        implements CYGINT_IO_SERIAL_LINE_STATUS_HW

        description   "
            This option includes the serial device driver for the 
            Cerfpda port 1."

        cdl_option CYGDAT_IO_SERIAL_ARM_CERFPDA_SERIAL1_NAME {
            display       "Device name for cerfpda serial port 1 driver"
            flavor        data
            default_value {"\"/dev/ser1\""}
            description   "
                This option specifies the name of the serial device
                for the Cerfpda port 1."
        }

        cdl_option CYGNUM_IO_SERIAL_ARM_CERFPDA_SERIAL1_BAUD {
            display       "Baud rate for the cerfpda serial port 1 driver"
            flavor        data
            legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400
                            3600 4800 7200 9600 14400 19200 38400
                            57600 115200 230400 }
            default_value 38400
            description   "
                This option specifies the default baud rate (speed)
                for the Cerfpda port 1."
         }

         cdl_option CYGNUM_IO_SERIAL_ARM_CERFPDA_SERIAL1_BUFSIZE {
             display       "Buffer size for the cerfpda serial port 1 driver"
             flavor        data
             legal_values  0 to 8192
             default_value 128
             description   "
                 This option specifies the size of the internal
                 buffers used for the cerfpda port 1."
         }
    }

}

# EOF ser_arm_cerfpda.cdl
