# ====================================================================
#
#      flash_phycore229x.cdl
#
#      FLASH memory - Hardware support on Phytec phyCORE LPC229x board
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002, 2008 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Uwe Kindler
# Original data:  gthomas
# Contributors:   gthomas
# Date:           2007-11-21
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_FLASH_PHYCORE229X {
    display       "phyCORE-LPC229x board FLASH memory support"
    description   "FLASH memory device support for Phytec phyCORE-LPC229x board"

    parent        CYGPKG_IO_FLASH
    active_if     CYGPKG_IO_FLASH
    requires      CYGPKG_HAL_ARM_LPC2XXX

    compile       -library=libextras.a flash_phycore229x.c

    # Arguably this should do in the generic package
    # but then there is a logic loop so you can never enable it.
    cdl_interface CYGINT_DEVS_FLASH_AMD_AM29XXXXX_REQUIRED {
        display   "Generic AMD AM29XXXXX driver required"
    }

    implements    CYGINT_DEVS_FLASH_AMD_AM29XXXXX_REQUIRED
    
    cdl_option CYGHWR_DEVS_FLASH_PHYCORE229X_AM29DL800 {
        display     "AMD AM29DL800 device fitted"
        flavor      bool
        active_if   { CYGHWR_HAL_ARM_PHYCORE229X_FLASH == "AM29DL800" }
        requires    CYGHWR_DEVS_FLASH_AMD_AM29DL800
        calculated  { CYGHWR_HAL_ARM_PHYCORE229X_FLASH == "AM29DL800" ? 1 : 0 }
    }
    
    cdl_option CYGHWR_DEVS_FLASH_PHYCORE229X_AM29LV800 {
        display     "AMD AM29LV800 device fitted"
        flavor      bool
        active_if   { CYGHWR_HAL_ARM_PHYCORE229X_FLASH == "AM29LV800" }
        requires    CYGHWR_DEVS_FLASH_AMD_AM29LV800
        calculated  { CYGHWR_HAL_ARM_PHYCORE229X_FLASH == "AM29LV800" ? 1 : 0 }
    }
    
    cdl_option CYGHWR_DEVS_FLASH_PHYCORE229X_AM29LV160 {
        display     "AMD AM29LV160 device fitted"
        flavor      bool
        active_if   { CYGHWR_HAL_ARM_PHYCORE229X_FLASH == "AM29LV160" }
        requires    CYGHWR_DEVS_FLASH_AMD_AM29LV160
        calculated  { CYGHWR_HAL_ARM_PHYCORE229X_FLASH == "AM29LV160" ? 1 : 0 }
    }
    
    cdl_option CYGHWR_DEVS_FLASH_PHYCORE229X_AM29LV320 {
        display     "AMD AM29LV320 device fitted"
        flavor      bool
        active_if   { CYGHWR_HAL_ARM_PHYCORE229X_FLASH == "AM29LV320" }
        requires    CYGHWR_DEVS_FLASH_AMD_AM29LV320D
        calculated  { CYGHWR_HAL_ARM_PHYCORE229X_FLASH == "AM29LV320" ? 1 : 0 }
    }
}

# EOF flash_phycore229x.cdl
