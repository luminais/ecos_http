# ====================================================================
#
#      flash_asb2303.cdl
#
#      FLASH memory - Hardware support on Matsushita ASB2303
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      msalter
# Original data:  dhowells
# Contributors:
# Date:           2002-11-08
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_FLASH_MN10300_ASB2303 {
    display       "Matsushita MN10300 ASB2303 FLASH memory support"

    parent        CYGPKG_IO_FLASH
    active_if     CYGPKG_IO_FLASH
    requires      CYGPKG_HAL_MN10300_AM33_ASB

    compile       mn10300_asb2303_flash.c

    # Arguably this should do in the generic package
    # but then there is a logic loop so you can never enable it.
    cdl_interface CYGINT_DEVS_FLASH_AMD_AM29XXXXX_REQUIRED {
        display   "Generic AMD AM29XXXXX driver required"
    }

    cdl_option CYGHWR_DEVS_FLASH_MN10300_ASB2303_BANK {
        display       "Which flash bank to program"
        flavor        data
        legal_values  { "BootPROM" "SysFlash" }
        default_value { "SysFlash" }
        description   "
           This option controls which bank of flash will be programmable."
    }

    implements    CYGINT_DEVS_FLASH_AMD_AM29XXXXX_REQUIRED
    requires      CYGHWR_DEVS_FLASH_AMD_AM29DL322D
    requires      CYGHWR_DEVS_FLASH_AMD_AM29DL324D
    requires      CYGHWR_DEVS_FLASH_AMD_AM29LV800
}
