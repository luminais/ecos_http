# ====================================================================
#
#      spi_at91.cdl
#
#      Atmel AT91 (ARM) SPI driver configuration data 
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002, 2009 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Savin Zlobec <savin@elatec.si> 
# Date:           2004-08-25
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_SPI_ARM_AT91 {
    parent        CYGPKG_IO_SPI
    active_if     CYGPKG_IO_SPI
    display       "Atmel AT91 SPI driver"
    requires      CYGPKG_HAL_ARM_AT91
    requires      CYGPKG_ERROR
    hardware
    include_dir   cyg/io
    compile       spi_at91.c
    compile       -library=libextras.a spi_at91_init.cxx

    cdl_option CYGHWR_DEVS_SPI_ARM_AT91_BUS0 {
        display       "Enable support for SPI bus 0"
        flavor        bool
        default_value 1
        description   "Enable this option to add support for the first 
	               SPI peripheral. The most AT91 devices only have one bus" 
    }

    cdl_interface CYGINT_DEVS_SPI_ARM_AT91_HAS_BUS1 {
        description   "
            This interface is implemented by HALs for devices which have
            the second SPI bus controller."
    }
        

    cdl_option CYGHWR_DEVS_SPI_ARM_AT91_BUS1 {
	active_if     CYGINT_DEVS_SPI_ARM_AT_HAS_BUS1
        display       "Enable support for SPI bus 1"
        flavor        bool
        default_value 0
        description   "Enable this option to add support for the second 
	               SPI peripheral. The most AT91 devices only have one bus" 
    }

    cdl_component CYGPKG_DEVS_SPI_ARM_AT91_BUS0_CFG {
        active_if   CYGHWR_DEVS_SPI_ARM_AT91_BUS0
	display     "Configuration options for SPI Bus 0"
	flavor      none
	description "This is the configuration options for SPI Bus 0"
	
        cdl_option CYGHWR_DEVS_SPI_ARM_AT91_BUS0_PCSDEC {
            display       "Support 4 to 16 decoder of chip select signals."
            flavor        bool
            default_value 0
            description   "Enable this option if SPI peripheral chip 
                selects are connected through an 4 to 16 decoder."
        }

        cdl_option CYGDAT_DEVS_SPI_ARM_AT91_BUS0_NPCS0 {
            display       "PIO-Pin used for NPSC0"
            flavor        data
            default_value  {"AT91_SPI_NPCS0"}
            description   "Any GPIO pin is able to be used as the SPI driver
	                   uses GPIO to control the chip selects. Specify the pin
			   as \"AT91_GPIO_PA13\" or \"AT91_GPIO_PB5\" etc. Specify 
			   \"NONE\" if this chip select is to be disabled"
        }
	
        cdl_option CYGDAT_DEVS_SPI_ARM_AT91_BUS0_NPCS1 {
            display       "PIO-Pin used for NPSC1"
            flavor        data
            default_value  {"AT91_SPI_NPCS1"}
            description   "Any GPIO pin is able to be used as the SPI driver
	                   uses GPIO to control the chip selects. Specify the pin
			   as \"AT91_GPIO_PA13\" or \"AT91_GPIO_PB5\" etc. Specify 
			   \"NONE\" if this chip select is to be disabled"
        }
        cdl_option CYGDAT_DEVS_SPI_ARM_AT91_BUS0_NPCS2 {
            display       "PIO-Pin used for NPSC2"
            flavor        data
            default_value  {"AT91_SPI_NPCS2"}
            description   "Any GPIO pin is able to be used as the SPI driver
	                   uses GPIO to control the chip selects. Specify the pin
			   as \"AT91_GPIO_PA13\" or \"AT91_GPIO_PB5\" etc. Specify 
			   \"NONE\" if this chip select is to be disabled"
        }
        cdl_option CYGDAT_DEVS_SPI_ARM_AT91_BUS0_NPCS3 {
            display       "PIO-Pin used for NPSC3"
            flavor        data
            default_value  {"AT91_SPI_NPCS3"}
            description   "Any GPIO pin is able to be used as the SPI driver
	                   uses GPIO to control the chip selects. Specify the pin
			   as \"AT91_GPIO_PA13\" or \"AT91_GPIO_PB5\" etc. Specify 
			   \"NONE\" if this chip select is to be disabled"
        }

    }

    cdl_component CYGPKG_DEVS_SPI_ARM_AT91_BUS1_CFG {
        active_if   CYGHWR_DEVS_SPI_ARM_AT91_BUS1
	display     "Configuration options for SPI Bus 1"
	flavor      none
	description "This is the configuration options for SPI Bus 1"
	
        cdl_option CYGHWR_DEVS_SPI_ARM_AT91_BUS1_PCSDEC {
            display       "Support 4 to 16 decoder of chip select signals."
            flavor        bool
            default_value 0
            description   "Enable this option if SPI peripheral chip 
                selects are connected through an 4 to 16 decoder."
        }

        cdl_option CYGDAT_DEVS_SPI_ARM_AT91_BUS1_NPCS0 {
            display       "PIO-Pin used for NPSC0"
            flavor        data
            default_value  {"AT91_SPI1_NPCS0"}
            description   "Any GPIO pin is able to be used as the SPI driver
	                   uses GPIO to control the chip selects. Specify the pin
			   as \"AT91_GPIO_PA13\" or \"AT91_GPIO_PB5\" etc. Specify 
			   \"NONE\" if this chip select is to be disabled"
        }
	
        cdl_option CYGDAT_DEVS_SPI_ARM_AT91_BUS1_NPCS1 {
            display       "PIO-Pin used for NPSC1"
            flavor        data
            default_value  {"AT91_SPI1_NPCS1"}
            description   "Any GPIO pin is able to be used as the SPI driver
	                   uses GPIO to control the chip selects. Specify the pin
			   as \"AT91_GPIO_PA13\" or \"AT91_GPIO_PB5\" etc. Specify 
			   \"NONE\" if this chip select is to be disabled"
        }
        cdl_option CYGDAT_DEVS_SPI_ARM_AT91_BUS1_NPCS2 {
            display       "PIO-Pin used for NPSC2"
            flavor        data
            default_value  {"AT91_SPI1_NPCS2"}
            description   "Any GPIO pin is able to be used as the SPI driver
	                   uses GPIO to control the chip selects. Specify the pin
			   as \"AT91_GPIO_PA13\" or \"AT91_GPIO_PB5\" etc. Specify 
			   \"NONE\" if this chip select is to be disabled"
        }
        cdl_option CYGDAT_DEVS_SPI_ARM_AT91_BUS1_NPCS3 {
            display       "PIO-Pin used for NPSC3"
            flavor        data
            default_value  {"AT91_SPI1_NPCS3"}
            description   "Any GPIO pin is able to be used as the SPI driver
	                   uses GPIO to control the chip selects. Specify the pin
			   as \"AT91_GPIO_PA13\" or \"AT91_GPIO_PB5\" etc. Specify 
			   \"NONE\" if this chip select is to be disabled"
        }

    }

    
    cdl_component CYGPKG_DEVS_SPI_ARM_AT91_OPTIONS {
        display "Atmel AT91 SPI driver build options"
        flavor  none
        description   "
	        Package specific build options including control over
	        compiler flags used only in building this package,
	        and details of which tests are built."

        cdl_option CYGPKG_DEVS_SPI_ARM_AT91_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the SPI device. These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_DEVS_SPI_ARM_AT91_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the SPI device. These flags are removed from
                the set of global flags if present."
        }
    }
}

# EOF spi_at91.cdl
