# ====================================================================
#
#      819x_switch_drivers.cdl
#
#      Ethernet drivers - support for RealTek 819x ethernet controller
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      David Hsu
# Contributors:
# Date:           2009-11-13
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package RTLPKG_DEVS_ETH_RLTK_819X_SWITCH {
    display       "RealTek 819x ethernet switch driver"
    description   "Ethernet switch driver for RTL819x."

    parent        CYGPKG_IO_ETH_DRIVERS
    active_if	  CYGPKG_IO_ETH_DRIVERS
    #active_if     CYGPKG_HAL_MIPS_RLX
	implements    CYGINT_IO_ETH_MULTICAST
    
    # FIXME: This really belongs in the RealTek_819x package ?
    cdl_interface RTLINT_DEVS_ETH_RLTK_819X_SWITCH_REQUIRED {
        display   "RealTek 819x ethernet switch driver required"
    }

    define_proc {
        puts $::cdl_system_header "/***** ethernet driver proc output start *****/"
        puts $::cdl_system_header "#define RTLDAT_DEVS_ETH_RLTK_819X_SWITCH_INL \"devs_eth_rltk_819x_switch.inl\""
        puts $::cdl_system_header "#define RTLDAT_DEVS_ETH_RLTK_819X_SWITCH_CFG <pkgconf/devs_eth_rltk_819x_switch.h>"
        puts $::cdl_system_header "/*****  ethernet driver proc output end  *****/"
    }

    cdl_component RTLPKG_DEVS_ETH_RLTK_819X_SWITCH_ETH0 {
        display       "Ethernet port 0 driver"
        flavor        bool
        default_value 1

        implements CYGHWR_NET_DRIVERS
        implements CYGHWR_NET_DRIVER_ETH0
        implements RTLINT_DEVS_ETH_RLTK_819X_SWITCH_REQUIRED

        cdl_option RTLDAT_DEVS_ETH_RLTK_819X_SWITCH_ETH0_NAME {
            display       "Device name for the ETH0 ethernet port 0 driver"
            flavor        data
            default_value {"\"eth0\""}
            description   "
                This option sets the name of the ethernet device for the
                RealTek 819x ethernet port 0."
        }
    }

    cdl_component RTLPKG_DEVS_ETH_RLTK_819X_SWITCH_ETH1 {
        display       "Ethernet port 1 driver"
        flavor        bool
        default_value { CYGPKG_REDBOOT ? 0 : 1 }

        implements CYGHWR_NET_DRIVERS
        implements CYGHWR_NET_DRIVER_ETH1
        implements RTLINT_DEVS_ETH_RLTK_819X_SWITCH_REQUIRED
        
	cdl_option RTLDAT_DEVS_ETH_RLTK_819X_SWITCH_ETH1_NAME {
            display       "Device name for the ETH1 ethernet port 1 driver"
            flavor        data
            default_value {"\"eth1\""}
            description   "
                This option sets the name of the ethernet device for the
                RealTek 819x ethernet port 1."
        }

	cdl_option RTLPKG_DEVS_ETH_RLTK_819X_SWITCH_ETH1_BRIDGED {
            display "eth1 bridged"
            default_value 0
            description   ""
	}
    }

 cdl_component RTLPKG_DEVS_ETH_RLTK_819X_SWITCH_ETH2 {
        display       "Ethernet port 2 driver"
        flavor        bool
        default_value 1

        implements CYGHWR_NET_DRIVERS
        implements CYGHWR_NET_DRIVER_ETH2
        implements RTLINT_DEVS_ETH_RLTK_819X_SWITCH_REQUIRED

        cdl_option RTLDAT_DEVS_ETH_RLTK_819X_SWITCH_ETH2_NAME {
            display       "Device name for the ETH2 ethernet port 2 driver"
            flavor        data
            default_value {"\"eth2\""}
            description   "
                This option sets the name of the ethernet device for the
                RealTek 819x ethernet port 2."
        }
    }

   cdl_component RTLPKG_DEVS_ETH_RLTK_819X_SWITCH_ETH3 {
        display       "Ethernet port 3 driver"
        flavor        bool
        default_value 1

        implements CYGHWR_NET_DRIVERS
        implements CYGHWR_NET_DRIVER_ETH3
        implements RTLINT_DEVS_ETH_RLTK_819X_SWITCH_REQUIRED

        cdl_option RTLDAT_DEVS_ETH_RLTK_819X_SWITCH_ETH3_NAME {
            display       "Device name for the ETH3 ethernet port 3 driver"
            flavor        data
            default_value {"\"eth3\""}
            description   "
                This option sets the name of the ethernet device for the
                RealTek 819x ethernet port 3."
        }
    }

   cdl_component RTLPKG_DEVS_ETH_RLTK_819X_SWITCH_ETH4 {
        display       "Ethernet port 4 driver"
        flavor        bool
        default_value 1

        implements CYGHWR_NET_DRIVERS
        implements CYGHWR_NET_DRIVER_ETH4
        implements RTLINT_DEVS_ETH_RLTK_819X_SWITCH_REQUIRED

        cdl_option RTLDAT_DEVS_ETH_RLTK_819X_SWITCH_ETH4_NAME {
            display       "Device name for the ETH4 ethernet port 4 driver"
            flavor        data
            default_value {"\"eth4\""}
            description   "
                This option sets the name of the ethernet device for the
                RealTek 819x ethernet port 4."
        }
    }

    cdl_component RTLPKG_DEVS_ETH_RLTK_819X_SWITCH_ETH7 {
        display       "Ethernet virtual port 7 driver for bridge vlan"
        flavor        bool
        default_value 1
 
        implements CYGHWR_NET_DRIVERS
        implements CYGHWR_NET_DRIVER_ETH7
        implements RTLINT_DEVS_ETH_RLTK_819X_SWITCH_REQUIRED
 
        cdl_option RTLDAT_DEVS_ETH_RLTK_819X_SWITCH_ETH7_NAME {
            display       "Device name for the ETH7 ethernet virtual port 7 driver"
            flavor        data
            default_value {"\"eth7\""}
            description   "
                This option sets the name of the ethernet device for the
                RealTek 819x ethernet virtual port 7."
        }
    }

   cdl_component RTLPKG_DEVS_ETH_RLTK_819X_SWITCH_PETH0 {
        display       "Ethernet peth0"
        flavor        bool
        default_value 0
		define -file system.h CONFIG_RTL_CUSTOM_PASSTHRU
        implements CYGHWR_NET_DRIVERS
        implements CYGHWR_NET_DRIVER_ETH5
        implements RTLINT_DEVS_ETH_RLTK_819X_SWITCH_REQUIRED

        cdl_option RTLDAT_DEVS_ETH_RLTK_819X_SWITCH_PETH0_NAME {
            display       "Device name for the peth0 driver"
            flavor        data
            default_value {"\"peth0\""}
            description   "
                This option sets the name of the ethernet device for the
                RealTek 819x peth0."
        }
    } 
   # SNMP demands to know stuff; this sadly makes us break the neat
    # abstraction of the device having nothing exported.
    # include_files include/819x_info.h
    # and tell them that it is available
    define_proc {
	    puts $::cdl_system_header \
      "#define CYGBLD_DEVS_ETH_DEVICE_H <pkgconf/devs_eth_rltk_819x_switch.h>"

      puts $::cdl_header "#include RTLDAT_DEVS_ETH_RLTK_819X_SWITCH_CFG";
    }

    cdl_option RTLPKG_DEVS_ETH_RLTK_819X_HAVE_ETH {
      display "Have ethernet devices"
      active_if { RTLPKG_DEVS_ETH_RLTK_819X_SWITCH_ETH0 || RTLPKG_DEVS_ETH_RLTK_819X_SWITCH_ETH1 }
      description   ""
      compile -library=libextras.a if_819x.c eth865x.c swCore.c swNic_poll.c swTable.c vlanTable.c  rtl865x_igmpsnooping_new.c rtl865x_igmpsnooping_glue.c common/rtl865x_eventMgr.c rtl819x_swNic.c common/rtl865x_netif.c l2Driver/rtl865x_fdb.c rtl819x_swNic.c

	define -file system.h CONFIG_RTL_819X_SWCORE 
	define -file system.h CONFIG_RTL_LAYERED_DRIVER
	define -file system.h CONFIG_RTL_LAYERED_DRIVER_L2
      calculated { RTLPKG_DEVS_ETH_RLTK_819X_SWITCH_ETH0 || RTLPKG_DEVS_ETH_RLTK_819X_SWITCH_ETH1 }
    }

    cdl_option RTLDBG_DEVS_ETH_RLTK_819X_SWITCH_CHATTER {
      display "Print debugging messages"
      default_value 0
      description   "
        If this option is set, a lot of debugging messages are printed
        to the console to help debug the driver."
    }

	cdl_option RTLPKG_DEVS_ETH_RLTK_HW_NAT {
        display "support hw nat"
                flavor   bool
                default_value 0
                description ""
				compile -library=libextras.a l4Driver/rtl865x_asicL4.c l4Driver/rtl865x_nat.c                

				define -file system.h CONFIG_RTL_LAYERED_DRIVER_L4
				define -file system.h CONFIG_RTL_HARDWARE_NAT
         }

	cdl_option RTLPKG_DEVS_ETH_RLTK_HW_COMMON {
        display "support hw nat||hw multicast"
                flavor   bool
                default_value 0
                description ""
                compile -library=libextras.a l3Driver/rtl865x_ppp.c  l3Driver/rtl865x_arp.c l3Driver/rtl865x_route.c l3Driver/rtl865x_ip.c l3Driver/rtl865x_nexthop.c

                define -file system.h CONFIG_RTL_LAYERED_DRIVER_L3
               
         }

	cdl_option RTLPKG_DEVS_ETH_RLTK_EXCHANGE_PORTMASK {
        display "support exchange portmask"
                flavor   bool
                default_value 0
                description ""
                define -file system.h CONFIG_RTL_EXCHANGE_PORTMASK
         }

	cdl_option RTLPKG_DEVS_ETH_RLTK_8367R {
        display "support 8367r"
                flavor   bool
                default_value 0
                description ""
                compile -library=libextras.a rtl8367r/rtk_api.c rtl8367r/rtl8367b_asicdrv_acl.c rtl8367r/rtl8367b_asicdrv.c rtl8367r/rtl8367b_asicdrv_cputag.c rtl8367r/rtl8367b_asicdrv_dot1x.c rtl8367r/rtl8367b_asicdrv_eav.c rtl8367r/rtl8367b_asicdrv_eee.c rtl8367r/rtl8367b_asicdrv_fc.c rtl8367r/rtl8367b_asicdrv_green.c rtl8367r/rtl8367b_asicdrv_hsb.c rtl8367r/rtl8367b_asicdrv_igmp.c rtl8367r/rtl8367b_asicdrv_inbwctrl.c rtl8367r/rtl8367b_asicdrv_interrupt.c rtl8367r/rtl8367b_asicdrv_led.c rtl8367r/rtl8367b_asicdrv_lut.c rtl8367r/rtl8367b_asicdrv_meter.c rtl8367r/rtl8367b_asicdrv_mib.c rtl8367r/rtl8367b_asicdrv_mirror.c rtl8367r/rtl8367b_asicdrv_misc.c rtl8367r/rtl8367b_asicdrv_phy.c rtl8367r/rtl8367b_asicdrv_port.c rtl8367r/rtl8367b_asicdrv_portIsolation.c rtl8367r/rtl8367b_asicdrv_qos.c rtl8367r/rtl8367b_asicdrv_rma.c rtl8367r/rtl8367b_asicdrv_scheduling.c rtl8367r/rtl8367b_asicdrv_storm.c rtl8367r/rtl8367b_asicdrv_svlan.c rtl8367r/rtl8367b_asicdrv_trunking.c rtl8367r/rtl8367b_asicdrv_unknownMulticast.c rtl8367r/rtl8367b_asicdrv_vlan.c common/gpio.c common/smi.c
                
				define -file system.h CONFIG_RTL_8367R_SUPPORT
         }

	cdl_option RTLPKG_DEVS_ETH_RLTK_8211E {
	display "support 8211E"
		flavor   bool
		default_value 0
		description ""
		define -file system.h CONFIG_RTL_8211E_SUPPORT
         }

	cdl_option RTLPKG_DEVS_ETH_RLTK_8211F {
       	display "support 8211F"
                flavor   bool
                default_value 0
                description ""
                define -file system.h CONFIG_RTL_8211F_SUPPORT
         }
	
	cdl_option RTLPKG_DEVS_ULINKER {
	        display "support ulinker"
                flavor   bool
                default_value 0
                description ""
                define -file system.h CONFIG_RTL_ULINKER
         }

	cdl_option RTLPKG_DEVS_ETH_RLTK_865x_IGMPSNOOPING {
    	display "support igmp snooping"
		flavor   bool
		default_value 0
		description ""
		#compile \
		#	rtl865x_igmpsnooping_new.c rtl865x_igmpsnooping_glue.c
		define -file system.h CONFIG_RTL_IGMP_SNOOPING
	 }


	cdl_option RTLPKG_DEVS_ETH_RLTK_865x_MLDSNOOPING {
        display "support mld snooping"
        flavor   bool
        default_value 0
        description ""
        define -file system.h CONFIG_RTL_MLD_SNOOPING
		active_if RTLPKG_DEVS_ETH_RLTK_865x_IGMPSNOOPING
     }
	
	cdl_option RTLPKG_DEVS_ETH_RLTK_865x_HW_MULTICAST {
		display "support hardware multicast"
		flavor bool
		default_value 0
		description ""
		compile -library=libextras.a rtl865x_multicast.c
		define -file system.h CONFIG_RTL_HARDWARE_MULTICAST
	}

        cdl_option RTLPKG_DEVS_ETH_RLTK_865x_PHYPOWERCTRL {
        display "support phy power on/off control"
        flavor   bool
        default_value 0
        description ""
        define -file system.h CONFIG_RTL_PHY_POWER_CTRL
     }

    cdl_component RTLPKG_DEVS_ETH_RLTK_819X_SWITCH_OPTIONS {
        display "819x ethernet support build options"
        flavor  none
	no_define

        cdl_option RTLPKG_DEVS_ETH_RLTK_819X_SWITCH_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "-D_KERNEL -D__ECOS -include pkgconf/system.h" }
            description   "
                This option modifies the set of compiler flags for
                building the 819x ethernet support package. These flags are used in addition
                to the set of global flags."
        }
    }
}

