# ====================================================================
#
#      sh_se77x9_eth_drivers.cdl
#
#      Ethernet drivers - support for NS DP83902A ethernet controller
#      on the Hitachi SE77X9 board.
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Contributors:   jskov
# Date:           2001-06-13
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_ETH_SH_SE77X9 {
    display       "SH SE77X9 board ethernet driver"
    description   "Ethernet driver for SH SE77X9 board."

    parent        CYGPKG_IO_ETH_DRIVERS
    active_if	  CYGPKG_IO_ETH_DRIVERS
    active_if     CYGPKG_HAL_SH_SH77X9_SE77X9

    include_dir   cyg/io

    # FIXME: This really belongs in the NS DP83902A package
    cdl_interface CYGINT_DEVS_ETH_NS_DP83902A_REQUIRED {
        display   "NS DP83902A ethernet driver required"
    }

    define_proc {
        puts $::cdl_system_header "/***** ethernet driver proc output start *****/"
        puts $::cdl_system_header "#define CYGDAT_DEVS_ETH_NS_DP83902A_INL <cyg/io/devs_eth_sh_se77x9.inl>"
        puts $::cdl_system_header "#define CYGDAT_DEVS_ETH_NS_DP83902A_CFG <pkgconf/devs_eth_sh_se77x9.h>"
        puts $::cdl_system_header "/*****  ethernet driver proc output end  *****/"
    }

    cdl_component CYGPKG_DEVS_ETH_SH_SE77X9_ETH0 {
        display       "SE77X9 ethernet port driver"
        flavor        bool
        default_value 1
        description   "
            This option includes the ethernet device driver for the
            SE77X9 port."

        implements CYGINT_DEVS_ETH_NS_DP83902A_REQUIRED

        cdl_option CYGDAT_DEVS_ETH_SH_SE77X9_ETH0_NAME {
            display       "Device name for the ETH0 ethernet driver"
            flavor        data
            default_value {"\"eth0\""}
            description   "
                This option sets the name of the ethernet device."
        }

        cdl_component CYGSEM_DEVS_ETH_SH_SE77X9_ETH0_SET_ESA {
            display       "Set the ethernet station address"
            flavor        bool
            calculated    1
            description   "Enabling this option will allow the ethernet
            station address to be forced to the value set by the
            configuration.  This may be required if the hardware does
            not include a serial EEPROM for the ESA."
            
            cdl_option CYGDAT_DEVS_ETH_SH_SE77X9_ETH0_ESA {
                display       "The ethernet station address"
                flavor        data
                default_value {"{0x08, 0x88, 0x12, 0x34, 0x56, 0x78}"}
                description   "The ethernet station address"
            }
        }
    }
}
