# ====================================================================
#
#      flash_mpc50.cdl
#
#      MPC 5.0 flash package configuration data
#
# ====================================================================
# ####ECOSGPLCOPYRIGHTBEGIN####                                             
# -------------------------------------------                               
# This file is part of eCos, the Embedded Configurable Operating System.    
# Copyright (C) 1998, 1999, 2000, 2001, 2002 Free Software Foundation, Inc. 
#
# eCos is free software; you can redistribute it and/or modify it under     
# the terms of the GNU General Public License as published by the Free      
# Software Foundation; either version 2 or (at your option) any later       
# version.                                                                  
#
# eCos is distributed in the hope that it will be useful, but WITHOUT       
# ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or     
# FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License     
# for more details.                                                         
#
# You should have received a copy of the GNU General Public License         
# along with eCos; if not, write to the Free Software Foundation, Inc.,     
# 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.             
#
# As a special exception, if other files instantiate templates or use       
# macros or inline functions from this file, or you compile this file       
# and link it with other works to produce a work based on this file,        
# this file does not by itself cause the resulting work to be covered by    
# the GNU General Public License. However the source code for this file     
# must still be made available in accordance with section (3) of the GNU    
# General Public License v2.                                                
#
# This exception does not invalidate any other reasons why a work based     
# on this file might be covered by the GNU General Public License.          
# -------------------------------------------                               
# ####ECOSGPLCOPYRIGHTEND####                                               
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      woehler
# Date:           2002-09-02
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_FLASH_MPC50 {
	display       "MPC 5.0 FLASH memory support"
	description   "FLASH memory device support for MPC 5.0"

	parent        CYGPKG_IO_FLASH
	active_if	  CYGPKG_IO_FLASH
	requires	  CYGPKG_HAL_ARM_XSCALE_MPC50
	requires      CYGPKG_DEVS_FLASH_STRATA

	include_dir   cyg/io

	cdl_interface CYGINT_DEVS_FLASH_STRATA_REQUIRED {
		display   "Generic StrataFLASH driver required"
	}

	implements    CYGINT_DEVS_FLASH_STRATA_REQUIRED

	define_proc {
		puts $::cdl_system_header "#define CYGDAT_DEVS_FLASH_STRATA_INL <cyg/io/mpc50_strataflash.inl>"
		puts $::cdl_system_header "#define CYGDAT_DEVS_FLASH_STRATA_CFG <pkgconf/devs_flash_mpc50.h>"
	}
}
