# ====================================================================
#
#      watchdog_sa11x0.cdl
#
#      eCos watchdog for ARM/SA11X0 driver configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Contributors:   hmt, jskov
# Date:           2001-02-27
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVICES_WATCHDOG_ARM_SA11X0 {
    parent        CYGPKG_IO_WATCHDOG
    active_if     CYGPKG_IO_WATCHDOG
    display       "SA11X0 watchdog driver"
    requires      CYGPKG_HAL_ARM_SA11X0
    requires      CYGPKG_KERNEL
    hardware
    compile       watchdog_sa11x0.cxx
    implements    CYGINT_WATCHDOG_HW_IMPLEMENTATIONS
    implements    CYGINT_WATCHDOG_RESETS_ON_TIMEOUT
    active_if     CYGIMP_WATCHDOG_HARDWARE

    cdl_option CYGIMP_WATCHDOG_HARDWARE {
        parent    CYGPKG_IO_WATCHDOG_IMPLEMENTATION
        display       "Hardware watchdog"
        default_value 1
        implements    CYGINT_WATCHDOG_IMPLEMENTATIONS
    }

    cdl_component CYGPKG_DEVICES_WATCHDOG_ARM_SA11X0_OPTIONS {
        display "SA11X0 watchdog build options"
        flavor  none
        description   "
	    Package specific build options including control over
	    compiler flags used only in building this package,
	    and details of which tests are built."


        cdl_option CYGPKG_DEVICES_WATCHDOG_ARM_SA11X0_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the watchdog device. These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_DEVICES_WATCHDOG_ARM_SA11X0_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the watchdog device. These flags are removed from
                the set of global flags if present."
        }

    }
}
