# ====================================================================
#
#      hal_arm_lpc2xxx_phycore229x.cdl
#
#      Phytec phyCORE-LPC2292/94 HAL package configuration data 
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002, 2008 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Uwe Kindler
# Contributors:   Uwe Kindler
# Date:           2007-11-20
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_ARM_LPC2XXX_PHYCORE229X {
    display       "Phytec phyCORE-LPC2292/94 development board HAL"
    parent        CYGPKG_HAL_ARM_LPC2XXX
    define_header hal_arm_lpc2xxx_phycore229x.h
    include_dir   cyg/hal
    hardware
    implements CYGINT_DEVS_CAN_LPC2XXX_CAN0
    implements CYGINT_DEVS_CAN_LPC2XXX_CAN1
    description   "
        The phyCORE-229x HAL package provides the support needed to run
        eCos on Phytec phyCORE-LPC2292/94 development board."

    compile       phycore229x_misc.c

    requires      { CYGHWR_HAL_ARM_LPC2XXX == "LPC2292" || CYGHWR_HAL_ARM_LPC2XXX == "LPC2294" }

    define_proc {
        puts $::cdl_system_header "#define CYGBLD_HAL_TARGET_H   <pkgconf/hal_arm.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_VARIANT_H  <pkgconf/hal_arm_lpc2xxx.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_PLATFORM_H <pkgconf/hal_arm_lpc2xxx_phycore229x.h>"
        puts $::cdl_header "#define HAL_PLATFORM_CPU    \"ARM7TDMI-S\""
        puts $::cdl_header "#define HAL_PLATFORM_BOARD  \"Phytec phyCORE-LPC2292/94\""
        puts $::cdl_header "#define HAL_PLATFORM_EXTRA  \"\""
    }

    cdl_component CYG_HAL_STARTUP {
        display       "Startup type"
        flavor        data
        default_value {"ROM"}
        legal_values  {"RAM" "ROM"}
        no_define
        define -file system.h CYG_HAL_STARTUP
        description   "
            Choose RAM or ROM startup type. Typically ROM startup is used for
            building RedBoot. RedBoot runs from internal on chip flash of
            LPC229x. Use RAM startup for building eCos applications.
            RedBoot manages the external on board flash devices. It copies
            the eCos application image from FLASH to phyCORE on board SRAM 
            and then starts the eCos application."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS {
        display      "Number of communication channels on the board"
        flavor       data
        calculated   2
        description "
            Channel 0: UART0, Channel 1: UART1"
    }
    
    
    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_DEFAULT {
        display      "Default console channel."
        active_if    CYGPRI_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_CONFIGURABLE
        flavor       data
        calculated   0
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL {
        display          "Debug serial port"
        active_if        CYGPRI_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_CONFIGURABLE
        flavor           data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        default_value    0
        description      "
            Phytec phyCORE-LPC2292/94 board has two serial channels. This option
            chooses which channel will be used to connect to a host
            running GDB."
     }

     cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL {
         display          "Diagnostic serial port"
         active_if        CYGPRI_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_CONFIGURABLE
         flavor data
         legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
         default_value    0
         description "
             The phyCORE-LPC2292/94 board has two serial ports. This option
             chooses which port will be used for diagnostic output."
     }

     cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_BAUD {
        display       "Diagnostic serial port baud rate"
        flavor        data
        legal_values  9600 19200 38400 57600 115200
        default_value 38400
        description   "
            This option selects the baud rate used for the diagnostic port."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_BAUD {
         display       "GDB serial port baud rate"
         flavor        data
         legal_values  9600 19200 38400 57600 115200
         default_value 38400
         description   "
             This option controls the baud rate used for the GDB
             connection."
    }
    
    cdl_component CYGHWR_HAL_ARM_PHYCORE229X_MEMCFG {
        display "Memory configuration"
        flavor  none
        description   "
            Configuration options for FLASH and SRAM memory of phyCORE
            board."
    
        cdl_option CYGHWR_HAL_ARM_PHYCORE229X_FLASH {
             display        "Flash configuration"
             flavor         data
             legal_values   { "AM29DL800" "AM29LV800" "AM29LV160" "AM29LV320" }
             default_value { "AM29LV800" }
             description    "
                 Select the type of FLASH device that is fitted on the phyCORE
                 board."       
        }
    
        cdl_option CYGHWR_HAL_ARM_PHYCORE229X_FLASH_DEVICE_SIZE {
            display       "FLASH device size"
            flavor        data
            calculated    { CYGHWR_HAL_ARM_PHYCORE229X_FLASH == "AM29DL800" ? 
                              0x100000 :
                            CYGHWR_HAL_ARM_PHYCORE229X_FLASH == "AM29LV800" ? 
                              0x100000 :
                            CYGHWR_HAL_ARM_PHYCORE229X_FLASH == "AM29LV160" ? 
                              0x200000 :
                            CYGHWR_HAL_ARM_PHYCORE229X_FLASH == "AM29LV320" ? 
                              0x400000 : 0x000 }
            description   "
                Size of one single flash device."                        
        }
    
        cdl_option CYGHWR_HAL_ARM_PHYCORE229X_FLASH_CNT {
            display        "Number of flash devices"
            flavor         data
            legal_values   { 0 2 4 }
            default_value  { 2 }
            description    "
                This option defines the number of flash devices
                fitted. The board supports two 16-bit data bus width
                Flash devices in parallel connected to a 32-bit data
                bus on the LPC2292/94. Flash devices are always fitted
                in pairs and there is space for up to 4 devices."
        }
    
        cdl_option CYGHWR_HAL_ARM_PHYCORE229X_FLASH_SIZE {
            display      "FLASH size"
            flavor        data
            calculated   { CYGHWR_HAL_ARM_PHYCORE229X_FLASH_DEVICE_SIZE * 
                           CYGHWR_HAL_ARM_PHYCORE229X_FLASH_CNT }
            description    "
                This option defines the size of the onboard FLASH. 
                The board can be fitted with 0, 2 or 4 FLASH devices of
                1MB, 2MB or 4MB."
        }
    
        cdl_option CYGHWR_HAL_ARM_PHYCORE229X_SRAM_SIZE {
            display       "SRAM size"
            flavor        data
            legal_values  { 0x100000 0x200000 0x400000 0x800000 }
            default_value 0x100000
            description   "
                This option defines the size of the onboard SRAM. 
                The board can be fittet with 2 or 4 SRAM devices of
                512KB, 1MB or 2MB."
        }
    }
    
    cdl_component CYGHWR_HAL_ARM_PHYCORE229X_ETH {
        display "Ethernet options"
        flavor  none
        description   "
            Configuration options for on board SMSC LAN91C111 ethernet 
            chip."
    
    
        cdl_option CYGHWR_HAL_ARM_PHYCORE229X_ETH_EINT {
            display       "Ethernet controller interrupt"
            flavor        data
            legal_values  { 0 1 }
            default_value { 0 }
            description   "
                Jumper J501 selects, which of the microcontroller external
                interrupts (EINT) connects with the interrupt output(LAN_IRQ) 
                of the Ethernet controller. This configuration option should 
                match the actual jumper settings. The LAN chip may use EINT0
                or EINT1."
        }
    
        cdl_option CYGHWR_HAL_ARM_PHYCORE229X_ETH_INT_PRIO {
            display       "Ethernet interrupt priority"
            flavor        data
            legal_values  { 0 to 16 }
            default_value { 15 }
            description   "
                Interrupt priority of ethernet interrupt.  The LPC2xxx
                eCos HAL supports up to 17 interrupt levels.
                Interrupt levels 0 - 15 are vectored IRQs. Vectored
                IRQs have a higher priority then non vectored IRQs and
                they are processed faster. Non vectored IRQs are all
                chained together into one single slot and the ISR need
                to find out which interrupt occured. The default value
                for the ethernt interrupt is 15.  This is the lowest
                vectored IRQ priority. That ensures that the ethernet
                interrupt is processed fast while it has still a lower
                priority than any other verctored interrupt."  
        }
    
        cdl_option CYGHWR_HAL_ARM_PHYCORE229X_ETH_MEM_AREA {
            display        "Ethernet controller memory area"
            flavor         data
            legal_values   { 0x82000000 0x83000000 }
            default_value  { 0x82000000 }
            description    "
                Access to the optional Ethernet controller can be established
                via /CS2 (addr. 0x82000000) or /CS3 (addr. 0x83000000) 
                configurable with Jumper J502. The default configuration 
                allows access via /CS2."
        }
    }

    # Real-time clock/counter specifics
    cdl_option CYGNUM_HAL_ARM_LPC2XXX_XTAL_FREQ {
        display       "CPU xtal frequency"
        flavor        data
        default_value {10000000}
    }

    cdl_option CYGNUM_HAL_ARM_LPC2XXX_PLL_MUL {
        display       "CPU PLL multiplier"
        flavor        data
        default_value {6}
    }

    cdl_option CYGNUM_HAL_ARM_LPC2XXX_CLOCK_SPEED {
        display       "CPU clock speed"
        flavor        data
        calculated { CYGNUM_HAL_ARM_LPC2XXX_PLL_MUL * 
                     CYGNUM_HAL_ARM_LPC2XXX_XTAL_FREQ }
    }
    
    cdl_component CYGBLD_GLOBAL_OPTIONS {
        display "Global build options"
        flavor  none
        parent  CYGPKG_NONE
        description   "
            Global build options including control over compiler flags,
            linker flags and choice of toolchain."

        cdl_option CYGBLD_GLOBAL_COMMAND_PREFIX {
            display "Global command prefix"
            flavor  data
            no_define
            default_value { "arm-eabi"}
            description "
                This option specifies the command prefix used when
                invoking the build tools."
        }

        cdl_option CYGBLD_GLOBAL_CFLAGS {
            display "Global compiler flags"
            flavor  data
            no_define
            default_value { CYGBLD_GLOBAL_WARNFLAGS . CYGBLD_ARCH_CFLAGS .
                            "-mcpu=arm7tdmi -g -O2 -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions " }
            description   "
                This option controls the global compiler flags which
                are used to compile all packages by default. Individual
                packages may define options which override these global
                flags."
        }

        cdl_option CYGBLD_GLOBAL_LDFLAGS {
            display "Global linker flags"
            flavor  data
            no_define
            default_value { CYGBLD_ARCH_LDFLAGS . "-mcpu=arm7tdmi -Wl,--gc-sections -Wl,-static -g -nostdlib" }
            description   "
                This option controls the global linker flags. Individual
                packages may define options which override these global
                flags."
        }
    }

    cdl_option CYGSEM_HAL_ROM_MONITOR {
        display       "Behave as a ROM monitor"
        flavor        bool
        default_value 0
        parent        CYGPKG_HAL_ROM_MONITOR
        requires      { CYG_HAL_STARTUP == "ROM"}
        description   "
            Enable this option if this program is to be used as a
            ROM monitor, i.e. applications will be loaded into RAM on
            the board, and this ROM monitor may process exceptions or
            interrupts generated from the application. This enables
            features such as utilizing a separate interrupt stack when
            exceptions are generated."
    }

    cdl_option CYGSEM_HAL_USE_ROM_MONITOR {
         display       "Work with a ROM monitor"
         flavor        booldata
         legal_values  { "Generic" "GDB_stubs" }
         default_value { CYG_HAL_STARTUP == "RAM" ? "GDB_stubs" : 0 }
         parent        CYGPKG_HAL_ROM_MONITOR
         requires      { CYG_HAL_STARTUP == "RAM" }
         description   "
             Support can be enabled for different varieties of ROM
             monitor.  This support changes various eCos semantics such
             as the encoding of diagnostic output, or the overriding of
             hardware interrupt vectors.
             Firstly there is \"Generic\" support which prevents the
             HAL from overriding the hardware vectors that it does not
             use, to instead allow an installed ROM monitor to handle
             them. This is the most basic support which is likely to be
             common to most implementations of ROM monitor.
             \"GDB_stubs\" provides support when GDB stubs are included
             in the ROM monitor or boot ROM."
    }

    cdl_component CYGPKG_REDBOOT_HAL_OPTIONS {
        display       "Redboot HAL options"
        flavor        none
        no_define
        parent        CYGPKG_REDBOOT
        active_if     CYGPKG_REDBOOT
        description   "
            This option lists the target's requirements for a valid
            Redboot configuration."

        cdl_option CYGBLD_BUILD_REDBOOT_BIN {
            display       "Build Redboot ROM binary image"
            active_if     CYGBLD_BUILD_REDBOOT
            requires      { !CYGBLD_BUILD_REDBOOT_WITH_EXEC }
            default_value 1
            no_define
            description "
                This option enables the conversion of the Redboot ELF
                image to a binary image suitable for ROM programming."

            make -priority 325 {
                <PREFIX>/bin/redboot.bin : <PREFIX>/bin/redboot.elf
                $(OBJCOPY) --strip-debug $< $(@:.bin=.img)
                $(OBJCOPY) -O srec $< $(@:.bin=.srec)
                $(OBJCOPY) -O ihex $< $(@:.bin=.hex)
                $(OBJCOPY) -O binary $< $@
            }

        }
    }

    cdl_component CYGHWR_MEMORY_LAYOUT {
        display "Memory layout"
        flavor data
        no_define
        calculated { (CYG_HAL_STARTUP == "RAM") ? "arm_lpc2xxx_phycore229x_ram" :
                                                  "arm_lpc2xxx_phycore229x_rom" }

        cdl_option CYGHWR_MEMORY_LAYOUT_LDI {
            display "Memory layout linker script fragment"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_LDI
            calculated { (CYG_HAL_STARTUP == "RAM") ? "<pkgconf/mlt_arm_lpc2xxx_phycore229x_ram.ldi>" :
                                                      "<pkgconf/mlt_arm_lpc2xxx_phycore229x_rom.ldi>" }
        }

        cdl_option CYGHWR_MEMORY_LAYOUT_H {
            display "Memory layout header file"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_H
            calculated { (CYG_HAL_STARTUP == "RAM") ? "<pkgconf/mlt_arm_lpc2xxx_phycore229x_ram.h>" :
                                                      "<pkgconf/mlt_arm_lpc2xxx_phycore229x_rom.h>" }
        }
    }
}
